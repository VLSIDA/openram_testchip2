VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO rram_test
  CLASS BLOCK ;
  FOREIGN rram_test ;
  ORIGIN 18.240 21.705 ;
  SIZE 65.120 BY 186.955 ;
  PIN p1T1R_WL
    ANTENNAGATEAREA 1.704000 ;
    PORT
      LAYER li1 ;
        RECT -4.520 1.505 -3.960 1.790 ;
        RECT -3.305 0.740 -2.745 1.025 ;
        RECT -2.255 -1.095 -1.695 -0.810 ;
        RECT -1.205 -5.105 -0.850 -4.820 ;
      LAYER mcon ;
        RECT -4.185 1.555 -4.015 1.725 ;
        RECT -2.970 0.790 -2.800 0.960 ;
        RECT -1.920 -1.045 -1.750 -0.875 ;
        RECT -1.115 -5.025 -0.945 -4.855 ;
      LAYER met1 ;
        RECT -4.320 1.025 -3.885 1.790 ;
        RECT -4.320 0.740 -2.670 1.025 ;
        RECT -4.320 -0.810 -3.885 0.740 ;
        RECT -4.320 -1.055 -1.620 -0.810 ;
        RECT -2.055 -4.655 -1.620 -1.055 ;
        RECT -2.055 -5.225 -0.695 -4.655 ;
      LAYER via ;
        RECT -4.235 1.530 -3.975 1.790 ;
        RECT -3.020 0.765 -2.760 1.025 ;
        RECT -1.970 -1.070 -1.710 -0.810 ;
        RECT -1.165 -5.065 -0.905 -4.805 ;
      LAYER met2 ;
        RECT -12.375 5.570 -10.560 7.350 ;
        RECT -11.010 1.790 -10.705 5.570 ;
        RECT -11.010 1.530 -3.885 1.790 ;
        RECT -3.105 0.765 -2.670 1.025 ;
        RECT -2.055 -1.070 -1.620 -0.810 ;
        RECT -1.350 -5.230 -0.690 -4.655 ;
    END
  END p1T1R_WL
  PIN p036_SL
    ANTENNADIFFAREA 0.108000 ;
    PORT
      LAYER li1 ;
        RECT -4.690 2.020 -4.520 2.350 ;
      LAYER mcon ;
        RECT -4.690 2.100 -4.520 2.270 ;
      LAYER met1 ;
        RECT -4.735 2.035 -4.415 2.355 ;
      LAYER via ;
        RECT -4.705 2.065 -4.445 2.325 ;
      LAYER met2 ;
        RECT -10.420 5.570 -8.605 7.350 ;
        RECT -9.110 2.355 -8.810 5.570 ;
        RECT -9.110 2.035 -4.415 2.355 ;
    END
  END p036_SL
  PIN p700_SL
    ANTENNADIFFAREA 2.100000 ;
    PORT
      LAYER li1 ;
        RECT -1.385 -3.000 -1.215 2.350 ;
      LAYER mcon ;
        RECT -1.385 1.965 -1.215 2.135 ;
        RECT -1.385 1.605 -1.215 1.775 ;
        RECT -1.385 1.245 -1.215 1.415 ;
        RECT -1.385 0.885 -1.215 1.055 ;
        RECT -1.385 0.525 -1.215 0.695 ;
        RECT -1.385 0.165 -1.215 0.335 ;
        RECT -1.385 -0.195 -1.215 -0.025 ;
        RECT -1.385 -0.555 -1.215 -0.385 ;
        RECT -1.385 -0.915 -1.215 -0.745 ;
        RECT -1.385 -1.275 -1.215 -1.105 ;
        RECT -1.385 -1.635 -1.215 -1.465 ;
        RECT -1.385 -1.995 -1.215 -1.825 ;
        RECT -1.385 -2.355 -1.215 -2.185 ;
        RECT -1.385 -2.715 -1.215 -2.545 ;
      LAYER met1 ;
        RECT -1.430 -3.000 -1.110 2.355 ;
      LAYER via ;
        RECT -1.400 1.890 -1.140 2.150 ;
        RECT -1.400 1.570 -1.140 1.830 ;
        RECT -1.400 1.250 -1.140 1.510 ;
        RECT -1.400 0.930 -1.140 1.190 ;
        RECT -1.400 0.610 -1.140 0.870 ;
        RECT -1.400 0.290 -1.140 0.550 ;
        RECT -1.400 -0.030 -1.140 0.230 ;
        RECT -1.400 -0.350 -1.140 -0.090 ;
        RECT -1.400 -0.670 -1.140 -0.410 ;
        RECT -1.400 -0.990 -1.140 -0.730 ;
        RECT -1.400 -1.310 -1.140 -1.050 ;
        RECT -1.400 -1.630 -1.140 -1.370 ;
        RECT -1.400 -1.950 -1.140 -1.690 ;
        RECT -1.400 -2.270 -1.140 -2.010 ;
        RECT -1.400 -2.590 -1.140 -2.330 ;
        RECT -1.400 -2.910 -1.140 -2.650 ;
      LAYER met2 ;
        RECT -18.240 5.570 -16.425 7.350 ;
        RECT -17.045 -2.310 -16.570 5.570 ;
        RECT -1.430 -2.310 -1.110 2.355 ;
        RECT -17.045 -2.600 -1.110 -2.310 ;
        RECT -1.430 -2.995 -1.110 -2.600 ;
    END
  END p700_SL
  PIN p300_SL
    ANTENNADIFFAREA 0.900000 ;
    PORT
      LAYER li1 ;
        RECT -2.420 -0.635 -2.250 2.350 ;
      LAYER mcon ;
        RECT -2.420 1.800 -2.250 1.970 ;
        RECT -2.420 1.440 -2.250 1.610 ;
        RECT -2.420 1.080 -2.250 1.250 ;
        RECT -2.420 0.720 -2.250 0.890 ;
        RECT -2.420 0.360 -2.250 0.530 ;
        RECT -2.420 0.000 -2.250 0.170 ;
        RECT -2.420 -0.360 -2.250 -0.190 ;
      LAYER met1 ;
        RECT -2.465 -0.635 -2.145 2.355 ;
      LAYER via ;
        RECT -2.435 1.810 -2.175 2.070 ;
        RECT -2.435 1.490 -2.175 1.750 ;
        RECT -2.435 1.170 -2.175 1.430 ;
        RECT -2.435 0.850 -2.175 1.110 ;
        RECT -2.435 0.530 -2.175 0.790 ;
        RECT -2.435 0.210 -2.175 0.470 ;
        RECT -2.435 -0.110 -2.175 0.150 ;
        RECT -2.435 -0.430 -2.175 -0.170 ;
      LAYER met2 ;
        RECT -16.285 5.570 -14.470 7.350 ;
        RECT -15.090 -0.175 -14.615 5.570 ;
        RECT -2.465 -0.175 -2.145 2.355 ;
        RECT -15.090 -0.435 -2.145 -0.175 ;
        RECT -2.465 -0.565 -2.145 -0.435 ;
    END
  END p300_SL
  PIN p100_SL
    ANTENNADIFFAREA 0.300000 ;
    PORT
      LAYER li1 ;
        RECT -3.475 1.400 -3.305 2.350 ;
      LAYER mcon ;
        RECT -3.475 1.980 -3.305 2.150 ;
        RECT -3.475 1.620 -3.305 1.790 ;
      LAYER met1 ;
        RECT -3.520 1.395 -3.200 2.355 ;
      LAYER via ;
        RECT -3.490 1.915 -3.230 2.175 ;
        RECT -3.490 1.595 -3.230 1.855 ;
      LAYER met2 ;
        RECT -14.330 5.570 -12.515 7.350 ;
        RECT -13.135 1.025 -12.760 5.570 ;
        RECT -3.520 1.360 -3.200 2.355 ;
        RECT -3.725 1.165 -3.200 1.360 ;
        RECT -3.725 1.025 -3.315 1.165 ;
        RECT -13.135 0.765 -3.520 1.025 ;
    END
  END p100_SL
  PIN RE_BR0
    ANTENNADIFFAREA 4.200000 ;
    PORT
      LAYER li1 ;
        RECT 18.825 -2.820 18.995 2.530 ;
        RECT 18.725 -19.420 18.895 -14.070 ;
      LAYER mcon ;
        RECT 18.825 2.145 18.995 2.315 ;
        RECT 18.825 1.785 18.995 1.955 ;
        RECT 18.825 1.425 18.995 1.595 ;
        RECT 18.825 1.065 18.995 1.235 ;
        RECT 18.825 0.705 18.995 0.875 ;
        RECT 18.825 0.345 18.995 0.515 ;
        RECT 18.825 -0.015 18.995 0.155 ;
        RECT 18.825 -0.375 18.995 -0.205 ;
        RECT 18.825 -0.735 18.995 -0.565 ;
        RECT 18.825 -1.095 18.995 -0.925 ;
        RECT 18.825 -1.455 18.995 -1.285 ;
        RECT 18.825 -1.815 18.995 -1.645 ;
        RECT 18.825 -2.175 18.995 -2.005 ;
        RECT 18.825 -2.535 18.995 -2.365 ;
        RECT 18.725 -14.455 18.895 -14.285 ;
        RECT 18.725 -14.815 18.895 -14.645 ;
        RECT 18.725 -15.175 18.895 -15.005 ;
        RECT 18.725 -15.535 18.895 -15.365 ;
        RECT 18.725 -15.895 18.895 -15.725 ;
        RECT 18.725 -16.255 18.895 -16.085 ;
        RECT 18.725 -16.615 18.895 -16.445 ;
        RECT 18.725 -16.975 18.895 -16.805 ;
        RECT 18.725 -17.335 18.895 -17.165 ;
        RECT 18.725 -17.695 18.895 -17.525 ;
        RECT 18.725 -18.055 18.895 -17.885 ;
        RECT 18.725 -18.415 18.895 -18.245 ;
        RECT 18.725 -18.775 18.895 -18.605 ;
        RECT 18.725 -19.135 18.895 -18.965 ;
      LAYER met1 ;
        RECT 18.780 -3.080 19.100 2.535 ;
        RECT 18.780 -3.285 21.695 -3.080 ;
        RECT 21.415 -4.970 21.695 -3.285 ;
        RECT 18.680 -19.680 19.000 -14.065 ;
        RECT 18.680 -19.885 21.595 -19.680 ;
        RECT 21.315 -21.570 21.595 -19.885 ;
      LAYER via ;
        RECT 18.810 2.070 19.070 2.330 ;
        RECT 18.810 1.750 19.070 2.010 ;
        RECT 18.810 1.430 19.070 1.690 ;
        RECT 18.810 1.110 19.070 1.370 ;
        RECT 18.810 0.790 19.070 1.050 ;
        RECT 18.810 0.470 19.070 0.730 ;
        RECT 18.810 0.150 19.070 0.410 ;
        RECT 18.810 -0.170 19.070 0.090 ;
        RECT 18.810 -0.490 19.070 -0.230 ;
        RECT 18.810 -0.810 19.070 -0.550 ;
        RECT 18.810 -1.130 19.070 -0.870 ;
        RECT 18.810 -1.450 19.070 -1.190 ;
        RECT 18.810 -1.770 19.070 -1.510 ;
        RECT 18.810 -2.090 19.070 -1.830 ;
        RECT 18.810 -2.410 19.070 -2.150 ;
        RECT 18.810 -2.730 19.070 -2.470 ;
        RECT 21.420 -4.910 21.680 -4.650 ;
        RECT 18.710 -14.530 18.970 -14.270 ;
        RECT 18.710 -14.850 18.970 -14.590 ;
        RECT 18.710 -15.170 18.970 -14.910 ;
        RECT 18.710 -15.490 18.970 -15.230 ;
        RECT 18.710 -15.810 18.970 -15.550 ;
        RECT 18.710 -16.130 18.970 -15.870 ;
        RECT 18.710 -16.450 18.970 -16.190 ;
        RECT 18.710 -16.770 18.970 -16.510 ;
        RECT 18.710 -17.090 18.970 -16.830 ;
        RECT 18.710 -17.410 18.970 -17.150 ;
        RECT 18.710 -17.730 18.970 -17.470 ;
        RECT 18.710 -18.050 18.970 -17.790 ;
        RECT 18.710 -18.370 18.970 -18.110 ;
        RECT 18.710 -18.690 18.970 -18.430 ;
        RECT 18.710 -19.010 18.970 -18.750 ;
        RECT 18.710 -19.330 18.970 -19.070 ;
        RECT 21.320 -21.510 21.580 -21.250 ;
      LAYER met2 ;
        RECT 19.175 8.070 20.990 9.850 ;
        RECT 20.660 5.220 20.990 8.070 ;
        RECT 20.660 4.990 21.700 5.220 ;
        RECT 18.780 -2.815 19.100 2.535 ;
        RECT 21.195 -4.580 21.700 4.990 ;
        RECT 18.680 -19.415 19.000 -14.065 ;
        RECT 21.190 -14.970 21.695 -4.580 ;
        RECT 21.185 -16.000 21.695 -14.970 ;
        RECT 21.190 -21.180 21.695 -16.000 ;
        RECT 21.090 -21.570 21.695 -21.180 ;
    END
  END RE_BR0
  PIN BL0
    ANTENNADIFFAREA 0.244800 ;
    PORT
      LAYER li1 ;
        RECT 16.165 0.530 17.505 0.780 ;
        RECT 16.065 -16.070 17.405 -15.820 ;
      LAYER mcon ;
        RECT 16.475 0.570 16.645 0.740 ;
        RECT 16.375 -16.030 16.545 -15.860 ;
      LAYER met1 ;
        RECT 15.855 2.845 16.695 3.405 ;
        RECT 16.435 0.780 16.695 2.845 ;
        RECT 16.415 0.510 16.705 0.780 ;
        RECT 12.885 -4.200 13.160 -3.980 ;
        RECT 16.435 -4.200 16.695 0.510 ;
        RECT 12.885 -4.405 16.695 -4.200 ;
        RECT 15.755 -13.755 16.595 -13.195 ;
        RECT 16.335 -15.820 16.595 -13.755 ;
        RECT 16.315 -16.090 16.605 -15.820 ;
        RECT 12.785 -20.800 13.060 -20.580 ;
        RECT 16.335 -20.800 16.595 -16.090 ;
        RECT 12.785 -21.005 16.595 -20.800 ;
      LAYER via ;
        RECT 16.015 3.000 16.275 3.260 ;
        RECT 12.890 -4.350 13.150 -4.090 ;
        RECT 15.915 -13.600 16.175 -13.340 ;
        RECT 12.790 -20.950 13.050 -20.690 ;
      LAYER met2 ;
        RECT 11.355 8.070 13.170 9.850 ;
        RECT 12.880 -20.575 13.170 8.070 ;
        RECT 15.855 3.400 16.425 3.410 ;
        RECT 15.030 3.120 16.425 3.400 ;
        RECT 15.855 2.835 16.425 3.120 ;
        RECT 15.755 -13.200 16.325 -13.190 ;
        RECT 14.930 -13.480 16.325 -13.200 ;
        RECT 15.755 -13.765 16.325 -13.480 ;
        RECT 12.780 -21.000 13.170 -20.575 ;
    END
  END BL0
  PIN RE_BL0
    ANTENNADIFFAREA 4.200000 ;
    PORT
      LAYER li1 ;
        RECT 14.550 -2.820 14.720 2.530 ;
        RECT 14.450 -19.420 14.620 -14.070 ;
      LAYER mcon ;
        RECT 14.550 2.145 14.720 2.315 ;
        RECT 14.550 1.785 14.720 1.955 ;
        RECT 14.550 1.425 14.720 1.595 ;
        RECT 14.550 1.065 14.720 1.235 ;
        RECT 14.550 0.705 14.720 0.875 ;
        RECT 14.550 0.345 14.720 0.515 ;
        RECT 14.550 -0.015 14.720 0.155 ;
        RECT 14.550 -0.375 14.720 -0.205 ;
        RECT 14.550 -0.735 14.720 -0.565 ;
        RECT 14.550 -1.095 14.720 -0.925 ;
        RECT 14.550 -1.455 14.720 -1.285 ;
        RECT 14.550 -1.815 14.720 -1.645 ;
        RECT 14.550 -2.175 14.720 -2.005 ;
        RECT 14.550 -2.535 14.720 -2.365 ;
        RECT 14.450 -14.455 14.620 -14.285 ;
        RECT 14.450 -14.815 14.620 -14.645 ;
        RECT 14.450 -15.175 14.620 -15.005 ;
        RECT 14.450 -15.535 14.620 -15.365 ;
        RECT 14.450 -15.895 14.620 -15.725 ;
        RECT 14.450 -16.255 14.620 -16.085 ;
        RECT 14.450 -16.615 14.620 -16.445 ;
        RECT 14.450 -16.975 14.620 -16.805 ;
        RECT 14.450 -17.335 14.620 -17.165 ;
        RECT 14.450 -17.695 14.620 -17.525 ;
        RECT 14.450 -18.055 14.620 -17.885 ;
        RECT 14.450 -18.415 14.620 -18.245 ;
        RECT 14.450 -18.775 14.620 -18.605 ;
        RECT 14.450 -19.135 14.620 -18.965 ;
      LAYER met1 ;
        RECT 14.505 -2.465 14.825 2.535 ;
        RECT 12.245 -2.780 14.825 -2.465 ;
        RECT 12.245 -4.925 12.610 -2.780 ;
        RECT 14.505 -2.820 14.825 -2.780 ;
        RECT 14.405 -19.065 14.725 -14.065 ;
        RECT 12.145 -19.380 14.725 -19.065 ;
        RECT 12.145 -21.525 12.510 -19.380 ;
        RECT 14.405 -19.420 14.725 -19.380 ;
      LAYER via ;
        RECT 14.535 2.070 14.795 2.330 ;
        RECT 14.535 1.750 14.795 2.010 ;
        RECT 14.535 1.430 14.795 1.690 ;
        RECT 14.535 1.110 14.795 1.370 ;
        RECT 14.535 0.790 14.795 1.050 ;
        RECT 14.535 0.470 14.795 0.730 ;
        RECT 14.535 0.150 14.795 0.410 ;
        RECT 14.535 -0.170 14.795 0.090 ;
        RECT 14.535 -0.490 14.795 -0.230 ;
        RECT 14.535 -0.810 14.795 -0.550 ;
        RECT 14.535 -1.130 14.795 -0.870 ;
        RECT 14.535 -1.450 14.795 -1.190 ;
        RECT 14.535 -1.770 14.795 -1.510 ;
        RECT 14.535 -2.090 14.795 -1.830 ;
        RECT 14.535 -2.410 14.795 -2.150 ;
        RECT 14.535 -2.730 14.795 -2.470 ;
        RECT 12.315 -4.910 12.575 -4.650 ;
        RECT 14.435 -14.530 14.695 -14.270 ;
        RECT 14.435 -14.850 14.695 -14.590 ;
        RECT 14.435 -15.170 14.695 -14.910 ;
        RECT 14.435 -15.490 14.695 -15.230 ;
        RECT 14.435 -15.810 14.695 -15.550 ;
        RECT 14.435 -16.130 14.695 -15.870 ;
        RECT 14.435 -16.450 14.695 -16.190 ;
        RECT 14.435 -16.770 14.695 -16.510 ;
        RECT 14.435 -17.090 14.695 -16.830 ;
        RECT 14.435 -17.410 14.695 -17.150 ;
        RECT 14.435 -17.730 14.695 -17.470 ;
        RECT 14.435 -18.050 14.695 -17.790 ;
        RECT 14.435 -18.370 14.695 -18.110 ;
        RECT 14.435 -18.690 14.695 -18.430 ;
        RECT 14.435 -19.010 14.695 -18.750 ;
        RECT 14.435 -19.330 14.695 -19.070 ;
        RECT 12.215 -21.510 12.475 -21.250 ;
      LAYER met2 ;
        RECT 9.400 8.070 11.215 9.850 ;
        RECT 10.900 5.220 11.215 8.070 ;
        RECT 10.900 4.865 12.740 5.220 ;
        RECT 12.235 -4.970 12.740 4.865 ;
        RECT 14.505 -2.815 14.825 2.535 ;
        RECT 12.235 -14.970 12.640 -4.970 ;
        RECT 12.235 -16.000 12.740 -14.970 ;
        RECT 12.235 -21.180 12.640 -16.000 ;
        RECT 14.405 -19.415 14.725 -14.065 ;
        RECT 12.135 -21.570 12.740 -21.180 ;
    END
  END RE_BL0
  PIN BR0
    ANTENNADIFFAREA 0.244800 ;
    PORT
      LAYER li1 ;
        RECT 16.165 -1.620 17.505 -1.370 ;
        RECT 16.065 -18.220 17.405 -17.970 ;
      LAYER mcon ;
        RECT 17.015 -1.580 17.185 -1.410 ;
        RECT 16.915 -18.180 17.085 -18.010 ;
      LAYER met1 ;
        RECT 16.955 2.840 17.845 3.420 ;
        RECT 16.955 0.780 17.245 2.840 ;
        RECT 16.965 -1.350 17.225 0.780 ;
        RECT 16.955 -1.620 17.245 -1.350 ;
        RECT 16.965 -4.200 17.225 -1.620 ;
        RECT 20.660 -4.200 20.935 -3.980 ;
        RECT 16.965 -4.405 20.935 -4.200 ;
        RECT 16.965 -4.410 17.225 -4.405 ;
        RECT 16.855 -13.760 17.745 -13.180 ;
        RECT 16.855 -15.820 17.145 -13.760 ;
        RECT 16.865 -17.950 17.125 -15.820 ;
        RECT 16.855 -18.220 17.145 -17.950 ;
        RECT 16.865 -20.800 17.125 -18.220 ;
        RECT 20.560 -20.800 20.835 -20.580 ;
        RECT 16.865 -21.005 20.835 -20.800 ;
        RECT 16.865 -21.010 17.125 -21.005 ;
      LAYER via ;
        RECT 17.425 2.990 17.685 3.250 ;
        RECT 20.665 -4.350 20.925 -4.090 ;
        RECT 17.325 -13.610 17.585 -13.350 ;
        RECT 20.565 -20.950 20.825 -20.690 ;
      LAYER met2 ;
        RECT 17.220 8.070 19.035 9.850 ;
        RECT 18.725 4.700 19.035 8.070 ;
        RECT 18.725 4.515 20.945 4.700 ;
        RECT 17.250 3.150 18.985 3.420 ;
        RECT 17.250 2.845 17.840 3.150 ;
        RECT 17.150 -13.450 18.885 -13.180 ;
        RECT 17.150 -13.755 17.740 -13.450 ;
        RECT 20.655 -20.575 20.945 4.515 ;
        RECT 20.555 -21.000 20.945 -20.575 ;
    END
  END BR0
  PIN p1T1R_TE
    PORT
      LAYER met2 ;
        RECT -8.465 5.570 -6.650 7.350 ;
        RECT -7.065 3.245 -6.650 5.570 ;
        RECT -7.065 3.240 -0.860 3.245 ;
        RECT -7.065 2.920 -4.530 3.240 ;
        RECT -4.210 2.920 -3.315 3.240 ;
        RECT -2.995 2.920 -2.260 3.240 ;
        RECT -1.940 2.920 -1.225 3.240 ;
        RECT -0.905 2.920 -0.860 3.240 ;
        RECT -7.065 2.900 -0.860 2.920 ;
    END
  END p1T1R_TE
  PIN p1R_SL
    PORT
      LAYER met1 ;
        RECT -5.710 4.435 -4.410 4.695 ;
      LAYER via ;
        RECT -5.670 4.435 -5.410 4.695 ;
      LAYER met2 ;
        RECT -6.510 5.570 -4.695 7.350 ;
        RECT -6.000 4.300 -5.055 5.570 ;
    END
  END p1R_SL
  PIN p1R_TE
    PORT
      LAYER met2 ;
        RECT -4.555 5.570 -2.740 7.350 ;
        RECT -4.555 4.725 -4.000 5.570 ;
        RECT -4.410 4.405 -4.000 4.725 ;
    END
  END p1R_TE
  PIN BR1
    ANTENNADIFFAREA 0.244800 ;
    PORT
      LAYER li1 ;
        RECT 36.415 -1.620 37.755 -1.370 ;
        RECT 36.315 -18.220 37.655 -17.970 ;
      LAYER mcon ;
        RECT 37.265 -1.580 37.435 -1.410 ;
        RECT 37.165 -18.180 37.335 -18.010 ;
      LAYER met1 ;
        RECT 37.205 2.840 38.095 3.420 ;
        RECT 37.205 0.780 37.495 2.840 ;
        RECT 37.215 -1.350 37.475 0.780 ;
        RECT 37.205 -1.620 37.495 -1.350 ;
        RECT 37.215 -4.200 37.475 -1.620 ;
        RECT 40.910 -4.200 41.185 -3.980 ;
        RECT 37.215 -4.405 41.185 -4.200 ;
        RECT 37.215 -4.410 37.475 -4.405 ;
        RECT 37.105 -13.760 37.995 -13.180 ;
        RECT 37.105 -15.820 37.395 -13.760 ;
        RECT 37.115 -17.950 37.375 -15.820 ;
        RECT 37.105 -18.220 37.395 -17.950 ;
        RECT 37.115 -20.800 37.375 -18.220 ;
        RECT 40.810 -20.800 41.085 -20.580 ;
        RECT 37.115 -21.005 41.085 -20.800 ;
        RECT 37.115 -21.010 37.375 -21.005 ;
      LAYER via ;
        RECT 37.675 2.990 37.935 3.250 ;
        RECT 40.915 -4.350 41.175 -4.090 ;
        RECT 37.575 -13.610 37.835 -13.350 ;
        RECT 40.815 -20.950 41.075 -20.690 ;
      LAYER met2 ;
        RECT 35.290 8.070 37.105 9.850 ;
        RECT 36.890 4.070 37.105 8.070 ;
        RECT 36.890 3.925 41.190 4.070 ;
        RECT 37.500 3.150 39.235 3.420 ;
        RECT 37.500 2.845 38.090 3.150 ;
        RECT 40.900 -3.975 41.190 3.925 ;
        RECT 37.400 -13.450 39.135 -13.180 ;
        RECT 37.400 -13.755 37.990 -13.450 ;
        RECT 40.905 -20.575 41.195 -3.975 ;
        RECT 40.805 -21.000 41.195 -20.575 ;
    END
  END BR1
  PIN RE_BR1
    ANTENNADIFFAREA 4.200000 ;
    PORT
      LAYER li1 ;
        RECT 39.075 -2.820 39.245 2.530 ;
        RECT 38.975 -19.420 39.145 -14.070 ;
      LAYER mcon ;
        RECT 39.075 2.145 39.245 2.315 ;
        RECT 39.075 1.785 39.245 1.955 ;
        RECT 39.075 1.425 39.245 1.595 ;
        RECT 39.075 1.065 39.245 1.235 ;
        RECT 39.075 0.705 39.245 0.875 ;
        RECT 39.075 0.345 39.245 0.515 ;
        RECT 39.075 -0.015 39.245 0.155 ;
        RECT 39.075 -0.375 39.245 -0.205 ;
        RECT 39.075 -0.735 39.245 -0.565 ;
        RECT 39.075 -1.095 39.245 -0.925 ;
        RECT 39.075 -1.455 39.245 -1.285 ;
        RECT 39.075 -1.815 39.245 -1.645 ;
        RECT 39.075 -2.175 39.245 -2.005 ;
        RECT 39.075 -2.535 39.245 -2.365 ;
        RECT 38.975 -14.455 39.145 -14.285 ;
        RECT 38.975 -14.815 39.145 -14.645 ;
        RECT 38.975 -15.175 39.145 -15.005 ;
        RECT 38.975 -15.535 39.145 -15.365 ;
        RECT 38.975 -15.895 39.145 -15.725 ;
        RECT 38.975 -16.255 39.145 -16.085 ;
        RECT 38.975 -16.615 39.145 -16.445 ;
        RECT 38.975 -16.975 39.145 -16.805 ;
        RECT 38.975 -17.335 39.145 -17.165 ;
        RECT 38.975 -17.695 39.145 -17.525 ;
        RECT 38.975 -18.055 39.145 -17.885 ;
        RECT 38.975 -18.415 39.145 -18.245 ;
        RECT 38.975 -18.775 39.145 -18.605 ;
        RECT 38.975 -19.135 39.145 -18.965 ;
      LAYER met1 ;
        RECT 39.030 -3.080 39.350 2.535 ;
        RECT 39.030 -3.285 41.945 -3.080 ;
        RECT 41.665 -4.970 41.945 -3.285 ;
        RECT 38.930 -19.680 39.250 -14.065 ;
        RECT 38.930 -19.885 41.845 -19.680 ;
        RECT 41.565 -21.570 41.845 -19.885 ;
      LAYER via ;
        RECT 39.060 2.070 39.320 2.330 ;
        RECT 39.060 1.750 39.320 2.010 ;
        RECT 39.060 1.430 39.320 1.690 ;
        RECT 39.060 1.110 39.320 1.370 ;
        RECT 39.060 0.790 39.320 1.050 ;
        RECT 39.060 0.470 39.320 0.730 ;
        RECT 39.060 0.150 39.320 0.410 ;
        RECT 39.060 -0.170 39.320 0.090 ;
        RECT 39.060 -0.490 39.320 -0.230 ;
        RECT 39.060 -0.810 39.320 -0.550 ;
        RECT 39.060 -1.130 39.320 -0.870 ;
        RECT 39.060 -1.450 39.320 -1.190 ;
        RECT 39.060 -1.770 39.320 -1.510 ;
        RECT 39.060 -2.090 39.320 -1.830 ;
        RECT 39.060 -2.410 39.320 -2.150 ;
        RECT 39.060 -2.730 39.320 -2.470 ;
        RECT 41.670 -4.910 41.930 -4.650 ;
        RECT 38.960 -14.530 39.220 -14.270 ;
        RECT 38.960 -14.850 39.220 -14.590 ;
        RECT 38.960 -15.170 39.220 -14.910 ;
        RECT 38.960 -15.490 39.220 -15.230 ;
        RECT 38.960 -15.810 39.220 -15.550 ;
        RECT 38.960 -16.130 39.220 -15.870 ;
        RECT 38.960 -16.450 39.220 -16.190 ;
        RECT 38.960 -16.770 39.220 -16.510 ;
        RECT 38.960 -17.090 39.220 -16.830 ;
        RECT 38.960 -17.410 39.220 -17.150 ;
        RECT 38.960 -17.730 39.220 -17.470 ;
        RECT 38.960 -18.050 39.220 -17.790 ;
        RECT 38.960 -18.370 39.220 -18.110 ;
        RECT 38.960 -18.690 39.220 -18.430 ;
        RECT 38.960 -19.010 39.220 -18.750 ;
        RECT 38.960 -19.330 39.220 -19.070 ;
        RECT 41.570 -21.510 41.830 -21.250 ;
      LAYER met2 ;
        RECT 37.245 8.070 39.060 9.850 ;
        RECT 38.795 4.395 39.060 8.070 ;
        RECT 38.795 4.210 41.945 4.395 ;
        RECT 39.030 -2.815 39.350 2.535 ;
        RECT 38.930 -19.415 39.250 -14.065 ;
        RECT 41.440 -14.970 41.945 4.210 ;
        RECT 41.435 -16.000 41.945 -14.970 ;
        RECT 41.440 -21.180 41.945 -16.000 ;
        RECT 41.340 -21.570 41.945 -21.180 ;
    END
  END RE_BR1
  PIN BL1
    ANTENNADIFFAREA 0.244800 ;
    PORT
      LAYER li1 ;
        RECT 36.415 0.530 37.755 0.780 ;
        RECT 36.315 -16.070 37.655 -15.820 ;
      LAYER mcon ;
        RECT 36.725 0.570 36.895 0.740 ;
        RECT 36.625 -16.030 36.795 -15.860 ;
      LAYER met1 ;
        RECT 36.105 2.845 36.945 3.405 ;
        RECT 36.685 0.780 36.945 2.845 ;
        RECT 36.665 0.510 36.955 0.780 ;
        RECT 33.135 -4.200 33.410 -3.980 ;
        RECT 36.685 -4.200 36.945 0.510 ;
        RECT 33.135 -4.405 36.945 -4.200 ;
        RECT 36.005 -13.755 36.845 -13.195 ;
        RECT 36.585 -15.820 36.845 -13.755 ;
        RECT 36.565 -16.090 36.855 -15.820 ;
        RECT 33.035 -20.800 33.310 -20.580 ;
        RECT 36.585 -20.800 36.845 -16.090 ;
        RECT 33.035 -21.005 36.845 -20.800 ;
      LAYER via ;
        RECT 36.265 3.000 36.525 3.260 ;
        RECT 33.140 -4.350 33.400 -4.090 ;
        RECT 36.165 -13.600 36.425 -13.340 ;
        RECT 33.040 -20.950 33.300 -20.690 ;
      LAYER met2 ;
        RECT 33.335 8.070 35.150 9.850 ;
        RECT 33.335 5.220 33.735 8.070 ;
        RECT 33.125 5.055 33.735 5.220 ;
        RECT 33.125 -3.975 33.415 5.055 ;
        RECT 36.105 3.400 36.675 3.410 ;
        RECT 35.280 3.120 36.675 3.400 ;
        RECT 36.105 2.835 36.675 3.120 ;
        RECT 33.130 -20.575 33.420 -3.975 ;
        RECT 36.005 -13.200 36.575 -13.190 ;
        RECT 35.180 -13.480 36.575 -13.200 ;
        RECT 36.005 -13.765 36.575 -13.480 ;
        RECT 33.030 -21.000 33.420 -20.575 ;
    END
  END BL1
  PIN RE_BL1
    ANTENNADIFFAREA 4.200000 ;
    PORT
      LAYER li1 ;
        RECT 34.800 -2.820 34.970 2.530 ;
        RECT 34.700 -19.420 34.870 -14.070 ;
      LAYER mcon ;
        RECT 34.800 2.145 34.970 2.315 ;
        RECT 34.800 1.785 34.970 1.955 ;
        RECT 34.800 1.425 34.970 1.595 ;
        RECT 34.800 1.065 34.970 1.235 ;
        RECT 34.800 0.705 34.970 0.875 ;
        RECT 34.800 0.345 34.970 0.515 ;
        RECT 34.800 -0.015 34.970 0.155 ;
        RECT 34.800 -0.375 34.970 -0.205 ;
        RECT 34.800 -0.735 34.970 -0.565 ;
        RECT 34.800 -1.095 34.970 -0.925 ;
        RECT 34.800 -1.455 34.970 -1.285 ;
        RECT 34.800 -1.815 34.970 -1.645 ;
        RECT 34.800 -2.175 34.970 -2.005 ;
        RECT 34.800 -2.535 34.970 -2.365 ;
        RECT 34.700 -14.455 34.870 -14.285 ;
        RECT 34.700 -14.815 34.870 -14.645 ;
        RECT 34.700 -15.175 34.870 -15.005 ;
        RECT 34.700 -15.535 34.870 -15.365 ;
        RECT 34.700 -15.895 34.870 -15.725 ;
        RECT 34.700 -16.255 34.870 -16.085 ;
        RECT 34.700 -16.615 34.870 -16.445 ;
        RECT 34.700 -16.975 34.870 -16.805 ;
        RECT 34.700 -17.335 34.870 -17.165 ;
        RECT 34.700 -17.695 34.870 -17.525 ;
        RECT 34.700 -18.055 34.870 -17.885 ;
        RECT 34.700 -18.415 34.870 -18.245 ;
        RECT 34.700 -18.775 34.870 -18.605 ;
        RECT 34.700 -19.135 34.870 -18.965 ;
      LAYER met1 ;
        RECT 34.755 -2.465 35.075 2.535 ;
        RECT 32.495 -2.780 35.075 -2.465 ;
        RECT 32.495 -4.925 32.860 -2.780 ;
        RECT 34.755 -2.820 35.075 -2.780 ;
        RECT 34.655 -19.065 34.975 -14.065 ;
        RECT 32.395 -19.380 34.975 -19.065 ;
        RECT 32.395 -21.525 32.760 -19.380 ;
        RECT 34.655 -19.420 34.975 -19.380 ;
      LAYER via ;
        RECT 34.785 2.070 35.045 2.330 ;
        RECT 34.785 1.750 35.045 2.010 ;
        RECT 34.785 1.430 35.045 1.690 ;
        RECT 34.785 1.110 35.045 1.370 ;
        RECT 34.785 0.790 35.045 1.050 ;
        RECT 34.785 0.470 35.045 0.730 ;
        RECT 34.785 0.150 35.045 0.410 ;
        RECT 34.785 -0.170 35.045 0.090 ;
        RECT 34.785 -0.490 35.045 -0.230 ;
        RECT 34.785 -0.810 35.045 -0.550 ;
        RECT 34.785 -1.130 35.045 -0.870 ;
        RECT 34.785 -1.450 35.045 -1.190 ;
        RECT 34.785 -1.770 35.045 -1.510 ;
        RECT 34.785 -2.090 35.045 -1.830 ;
        RECT 34.785 -2.410 35.045 -2.150 ;
        RECT 34.785 -2.730 35.045 -2.470 ;
        RECT 32.565 -4.910 32.825 -4.650 ;
        RECT 34.685 -14.530 34.945 -14.270 ;
        RECT 34.685 -14.850 34.945 -14.590 ;
        RECT 34.685 -15.170 34.945 -14.910 ;
        RECT 34.685 -15.490 34.945 -15.230 ;
        RECT 34.685 -15.810 34.945 -15.550 ;
        RECT 34.685 -16.130 34.945 -15.870 ;
        RECT 34.685 -16.450 34.945 -16.190 ;
        RECT 34.685 -16.770 34.945 -16.510 ;
        RECT 34.685 -17.090 34.945 -16.830 ;
        RECT 34.685 -17.410 34.945 -17.150 ;
        RECT 34.685 -17.730 34.945 -17.470 ;
        RECT 34.685 -18.050 34.945 -17.790 ;
        RECT 34.685 -18.370 34.945 -18.110 ;
        RECT 34.685 -18.690 34.945 -18.430 ;
        RECT 34.685 -19.010 34.945 -18.750 ;
        RECT 34.685 -19.330 34.945 -19.070 ;
        RECT 32.465 -21.510 32.725 -21.250 ;
      LAYER met2 ;
        RECT 31.180 8.070 32.995 9.850 ;
        RECT 32.480 -4.580 32.985 8.070 ;
        RECT 34.755 -2.815 35.075 2.535 ;
        RECT 32.485 -4.970 32.990 -4.580 ;
        RECT 32.485 -14.970 32.890 -4.970 ;
        RECT 32.485 -16.000 32.990 -14.970 ;
        RECT 32.485 -21.180 32.890 -16.000 ;
        RECT 34.655 -19.415 34.975 -14.065 ;
        RECT 32.385 -21.570 32.990 -21.180 ;
    END
  END RE_BL1
  PIN RE_WL1
    ANTENNAGATEAREA 4.200000 ;
    PORT
      LAYER li1 ;
        RECT 45.380 -20.675 45.780 -20.385 ;
        RECT 10.750 -20.845 22.820 -20.675 ;
        RECT 31.000 -20.845 45.780 -20.675 ;
        RECT 14.630 -21.525 14.985 -20.845 ;
        RECT 18.905 -21.525 19.260 -20.845 ;
        RECT 34.880 -21.525 35.235 -20.845 ;
        RECT 39.155 -21.525 39.510 -20.845 ;
      LAYER mcon ;
        RECT 22.565 -20.845 22.735 -20.675 ;
        RECT 31.110 -20.845 31.280 -20.675 ;
        RECT 45.485 -20.680 45.655 -20.510 ;
      LAYER met1 ;
        RECT 22.455 -20.995 31.365 -20.630 ;
        RECT 45.380 -20.805 45.780 -20.385 ;
      LAYER via ;
        RECT 45.455 -20.720 45.715 -20.460 ;
      LAYER met2 ;
        RECT 45.065 8.070 46.880 9.850 ;
        RECT 45.380 -20.845 45.780 8.070 ;
    END
  END RE_WL1
  PIN RE_WL0
    ANTENNAGATEAREA 4.200000 ;
    PORT
      LAYER li1 ;
        RECT 42.970 -4.075 43.370 -3.825 ;
        RECT 10.850 -4.245 22.725 -4.075 ;
        RECT 31.100 -4.245 45.870 -4.075 ;
        RECT 14.730 -4.925 15.085 -4.245 ;
        RECT 19.005 -4.925 19.360 -4.245 ;
        RECT 34.980 -4.925 35.335 -4.245 ;
        RECT 39.255 -4.925 39.610 -4.245 ;
      LAYER mcon ;
        RECT 22.470 -4.245 22.640 -4.075 ;
        RECT 31.210 -4.245 31.380 -4.075 ;
        RECT 43.075 -4.120 43.245 -3.950 ;
      LAYER met1 ;
        RECT 22.360 -4.395 31.465 -4.030 ;
        RECT 42.970 -4.245 43.370 -3.825 ;
      LAYER via ;
        RECT 43.045 -4.160 43.305 -3.900 ;
      LAYER met2 ;
        RECT 41.155 8.070 42.970 9.850 ;
        RECT 42.590 5.270 42.970 8.070 ;
        RECT 42.590 4.910 43.370 5.270 ;
        RECT 42.970 -4.245 43.370 4.910 ;
    END
  END RE_WL0
  PIN WL1
    ANTENNAGATEAREA 0.216000 ;
    PORT
      LAYER li1 ;
        RECT 15.290 -20.215 15.605 -19.660 ;
        RECT 35.540 -20.215 35.855 -19.660 ;
        RECT 43.820 -20.215 44.220 -19.925 ;
        RECT 10.750 -20.385 22.820 -20.215 ;
        RECT 31.000 -20.385 44.220 -20.215 ;
      LAYER mcon ;
        RECT 22.565 -20.385 22.735 -20.215 ;
        RECT 31.110 -20.385 31.280 -20.215 ;
        RECT 43.925 -20.220 44.095 -20.050 ;
      LAYER met1 ;
        RECT 22.455 -20.430 31.365 -20.040 ;
        RECT 43.820 -20.345 44.220 -19.925 ;
      LAYER via ;
        RECT 43.895 -20.260 44.155 -20.000 ;
      LAYER met2 ;
        RECT 43.110 8.070 44.925 9.850 ;
        RECT 43.820 -20.385 44.220 8.070 ;
    END
  END WL1
  PIN WL0
    ANTENNAGATEAREA 0.216000 ;
    PORT
      LAYER li1 ;
        RECT 15.390 -3.615 15.705 -3.060 ;
        RECT 35.640 -3.615 35.955 -3.060 ;
        RECT 42.270 -3.615 42.670 -3.365 ;
        RECT 10.850 -3.785 22.725 -3.615 ;
        RECT 31.100 -3.785 42.670 -3.615 ;
      LAYER mcon ;
        RECT 22.470 -3.785 22.640 -3.615 ;
        RECT 31.210 -3.785 31.380 -3.615 ;
        RECT 42.375 -3.660 42.545 -3.490 ;
      LAYER met1 ;
        RECT 22.360 -3.830 31.465 -3.440 ;
        RECT 42.270 -3.785 42.670 -3.365 ;
      LAYER via ;
        RECT 42.345 -3.700 42.605 -3.440 ;
      LAYER met2 ;
        RECT 39.200 8.070 41.015 9.850 ;
        RECT 40.605 4.695 41.010 8.070 ;
        RECT 40.605 4.535 42.670 4.695 ;
        RECT 42.270 -3.785 42.670 4.535 ;
    END
  END WL0
  PIN pVDD_HEADER0
    ANTENNAGATEAREA 0.108000 ;
    PORT
      LAYER li1 ;
        RECT 15.865 5.500 16.425 5.785 ;
        RECT 36.115 5.500 36.675 5.785 ;
      LAYER mcon ;
        RECT 16.200 5.565 16.370 5.735 ;
        RECT 36.450 5.565 36.620 5.735 ;
      LAYER met1 ;
        RECT 15.825 5.465 36.755 5.935 ;
      LAYER via ;
        RECT 23.375 5.555 23.635 5.815 ;
      LAYER met2 ;
        RECT 22.730 8.070 24.545 9.850 ;
        RECT 23.225 5.365 23.790 8.070 ;
    END
  END pVDD_HEADER0
  PIN pGND_HEADER0
    ANTENNAGATEAREA 0.108000 ;
    PORT
      LAYER li1 ;
        RECT 17.460 4.875 18.020 5.160 ;
        RECT 37.710 4.875 38.270 5.160 ;
      LAYER mcon ;
        RECT 17.795 4.940 17.965 5.110 ;
        RECT 38.045 4.940 38.215 5.110 ;
      LAYER met1 ;
        RECT 17.380 4.825 31.560 5.225 ;
        RECT 37.945 5.160 38.280 6.650 ;
        RECT 37.910 4.875 38.345 5.160 ;
      LAYER via ;
        RECT 37.985 6.355 38.245 6.615 ;
        RECT 25.500 4.885 25.760 5.145 ;
        RECT 31.180 4.900 31.440 5.160 ;
      LAYER met2 ;
        RECT 24.685 8.070 26.500 9.850 ;
        RECT 25.345 4.090 25.910 8.070 ;
        RECT 31.100 4.830 31.965 6.795 ;
        RECT 37.635 6.120 38.365 6.890 ;
      LAYER via2 ;
        RECT 31.370 6.385 31.650 6.665 ;
        RECT 37.970 6.345 38.250 6.625 ;
      LAYER met3 ;
        RECT 31.100 6.180 38.335 6.795 ;
    END
  END pGND_HEADER0
  PIN pVDD_HEADER1
    ANTENNAGATEAREA 0.108000 ;
    PORT
      LAYER li1 ;
        RECT 15.765 -11.100 16.325 -10.815 ;
        RECT 36.015 -11.100 36.575 -10.815 ;
      LAYER mcon ;
        RECT 16.100 -11.035 16.270 -10.865 ;
        RECT 36.350 -11.035 36.520 -10.865 ;
      LAYER met1 ;
        RECT 15.725 -10.815 36.425 -10.685 ;
        RECT 15.725 -11.100 36.650 -10.815 ;
        RECT 15.725 -11.155 36.425 -11.100 ;
      LAYER via ;
        RECT 27.775 -11.065 28.035 -10.805 ;
      LAYER met2 ;
        RECT 26.640 8.070 28.455 9.850 ;
        RECT 27.625 -11.255 28.190 8.070 ;
    END
  END pVDD_HEADER1
  PIN pGND_HEADER1
    ANTENNAGATEAREA 0.108000 ;
    PORT
      LAYER li1 ;
        RECT 17.360 -11.725 17.920 -11.440 ;
        RECT 37.610 -11.725 38.170 -11.440 ;
      LAYER mcon ;
        RECT 17.695 -11.660 17.865 -11.490 ;
        RECT 37.945 -11.660 38.115 -11.490 ;
      LAYER met1 ;
        RECT 37.710 -10.425 38.555 -9.660 ;
        RECT 17.280 -11.775 30.110 -11.375 ;
        RECT 37.810 -11.725 38.245 -10.425 ;
      LAYER via ;
        RECT 38.000 -10.175 38.260 -9.915 ;
        RECT 29.690 -11.700 29.950 -11.440 ;
      LAYER met2 ;
        RECT 28.595 8.070 30.410 9.850 ;
        RECT 29.545 -12.510 30.110 8.070 ;
        RECT 37.710 -10.425 38.555 -9.660 ;
      LAYER via2 ;
        RECT 29.685 -10.185 29.965 -9.905 ;
        RECT 37.985 -10.185 38.265 -9.905 ;
      LAYER met3 ;
        RECT 29.545 -10.250 38.435 -9.850 ;
    END
  END pGND_HEADER1
  PIN vccd1
    ANTENNADIFFAREA 1.132100 ;
    PORT
      LAYER nwell ;
        RECT 15.530 5.470 16.530 5.830 ;
        RECT 35.780 5.470 36.780 5.830 ;
        RECT 14.860 4.440 16.530 5.470 ;
        RECT 34.910 4.370 36.780 5.470 ;
        RECT 15.715 -2.505 16.695 0.780 ;
        RECT 35.965 -2.505 36.945 0.780 ;
        RECT 15.430 -11.130 16.430 -10.770 ;
        RECT 35.680 -11.130 36.680 -10.770 ;
        RECT 14.715 -12.075 16.430 -11.130 ;
        RECT 34.885 -12.245 36.680 -11.130 ;
        RECT 15.615 -19.105 16.595 -15.820 ;
        RECT 35.865 -19.105 36.845 -15.820 ;
      LAYER li1 ;
        RECT 14.950 4.940 15.865 5.270 ;
        RECT 35.265 4.940 36.115 5.270 ;
        RECT 15.915 -2.505 16.175 -1.925 ;
        RECT 36.165 -2.505 36.425 -1.925 ;
        RECT 14.840 -11.660 15.765 -11.330 ;
        RECT 35.010 -11.660 36.015 -11.330 ;
        RECT 15.815 -19.105 16.075 -18.525 ;
        RECT 36.065 -19.105 36.325 -18.525 ;
      LAYER mcon ;
        RECT 15.695 5.020 15.865 5.190 ;
        RECT 35.945 5.020 36.115 5.190 ;
        RECT 15.965 -2.360 16.135 -2.190 ;
        RECT 36.215 -2.360 36.385 -2.190 ;
        RECT 15.595 -11.580 15.765 -11.410 ;
        RECT 35.845 -11.580 36.015 -11.410 ;
        RECT 15.865 -18.960 16.035 -18.790 ;
        RECT 36.115 -18.960 36.285 -18.790 ;
      LAYER met1 ;
        RECT 13.440 6.710 35.115 7.135 ;
        RECT 14.840 4.935 15.970 5.255 ;
        RECT 35.260 4.935 36.220 5.255 ;
        RECT 13.440 -3.855 13.800 -3.685 ;
        RECT 15.915 -3.855 16.175 -2.035 ;
        RECT 13.440 -4.060 16.175 -3.855 ;
        RECT 33.690 -3.855 34.050 -3.685 ;
        RECT 36.165 -3.855 36.425 -2.035 ;
        RECT 33.690 -4.060 36.425 -3.855 ;
        RECT 14.820 -11.665 15.870 -11.345 ;
        RECT 34.935 -11.665 36.120 -11.345 ;
        RECT 13.340 -20.455 13.700 -20.285 ;
        RECT 15.815 -20.455 16.075 -18.635 ;
        RECT 13.340 -20.660 16.075 -20.455 ;
        RECT 33.590 -20.455 33.950 -20.285 ;
        RECT 36.065 -20.455 36.325 -18.635 ;
        RECT 33.590 -20.660 36.325 -20.455 ;
      LAYER via ;
        RECT 13.490 6.795 13.750 7.055 ;
        RECT 34.415 6.805 34.675 7.065 ;
        RECT 14.980 4.975 15.240 5.235 ;
        RECT 35.920 4.955 36.180 5.215 ;
        RECT 13.485 -3.995 13.745 -3.735 ;
        RECT 33.735 -3.995 33.995 -3.735 ;
        RECT 14.880 -11.625 15.140 -11.365 ;
        RECT 35.830 -11.645 36.090 -11.385 ;
        RECT 13.385 -20.595 13.645 -20.335 ;
        RECT 33.635 -20.595 33.895 -20.335 ;
      LAYER met2 ;
        RECT 13.435 8.075 15.250 9.855 ;
        RECT 13.440 -20.280 13.805 8.075 ;
        RECT 34.055 6.700 35.110 7.570 ;
        RECT 14.495 4.685 15.350 5.545 ;
        RECT 34.055 4.760 34.420 6.700 ;
        RECT 35.800 4.815 36.330 5.505 ;
        RECT 33.685 4.150 34.420 4.760 ;
        RECT 33.685 -3.680 34.055 4.150 ;
        RECT 14.395 -11.915 15.250 -11.055 ;
        RECT 33.690 -20.280 34.055 -3.680 ;
        RECT 35.460 -11.860 36.280 -11.235 ;
        RECT 13.340 -20.660 13.805 -20.280 ;
        RECT 33.590 -20.660 34.055 -20.280 ;
      LAYER via2 ;
        RECT 13.705 9.250 13.985 9.530 ;
        RECT 14.190 9.250 14.470 9.530 ;
        RECT 14.700 9.250 14.980 9.530 ;
        RECT 13.705 8.835 13.985 9.115 ;
        RECT 14.190 8.835 14.470 9.115 ;
        RECT 14.700 8.835 14.980 9.115 ;
        RECT 13.705 8.395 13.985 8.675 ;
        RECT 14.190 8.395 14.470 8.675 ;
        RECT 14.700 8.395 14.980 8.675 ;
        RECT 14.655 4.970 14.935 5.250 ;
        RECT 35.910 5.090 36.190 5.370 ;
        RECT 14.555 -11.630 14.835 -11.350 ;
        RECT 35.750 -11.735 36.030 -11.455 ;
      LAYER met3 ;
        RECT 13.435 8.075 15.250 9.855 ;
        RECT 14.495 5.465 15.350 5.545 ;
        RECT 14.495 4.975 36.275 5.465 ;
        RECT 14.495 4.685 15.350 4.975 ;
        RECT 14.395 -11.430 36.100 -11.055 ;
        RECT 14.395 -11.915 15.250 -11.430 ;
        RECT 35.680 -11.805 36.100 -11.430 ;
      LAYER via3 ;
        RECT 13.685 9.230 14.005 9.550 ;
        RECT 14.170 9.230 14.490 9.550 ;
        RECT 14.680 9.230 15.000 9.550 ;
        RECT 13.685 8.815 14.005 9.135 ;
        RECT 14.170 8.815 14.490 9.135 ;
        RECT 14.680 8.815 15.000 9.135 ;
        RECT 13.685 8.375 14.005 8.695 ;
        RECT 14.170 8.375 14.490 8.695 ;
        RECT 14.680 8.375 15.000 8.695 ;
        RECT 14.635 4.950 14.955 5.270 ;
        RECT 14.535 -11.650 14.855 -11.330 ;
      LAYER met4 ;
        RECT 13.435 -16.000 15.250 164.000 ;
    END
  END vccd1
  PIN vssd1
    ANTENNADIFFAREA 0.432000 ;
    PORT
      LAYER li1 ;
        RECT 17.290 4.315 17.460 4.645 ;
        RECT 37.540 4.315 37.710 4.645 ;
        RECT -6.145 3.565 -2.240 4.025 ;
        RECT -6.145 -1.395 -5.315 3.565 ;
        RECT -6.145 -2.230 -2.155 -1.395 ;
        RECT 17.490 -2.505 17.750 -1.925 ;
        RECT 37.740 -2.505 38.000 -1.925 ;
        RECT 17.190 -12.285 17.360 -11.955 ;
        RECT 37.440 -12.285 37.610 -11.955 ;
        RECT 17.390 -19.105 17.650 -18.525 ;
        RECT 37.640 -19.105 37.900 -18.525 ;
      LAYER mcon ;
        RECT 17.290 4.395 17.460 4.565 ;
        RECT 37.540 4.395 37.710 4.565 ;
        RECT -5.460 3.720 -5.290 3.890 ;
        RECT -4.990 3.715 -4.820 3.885 ;
        RECT -4.465 3.705 -4.295 3.875 ;
        RECT -3.995 3.700 -3.825 3.870 ;
        RECT -3.570 3.710 -3.400 3.880 ;
        RECT -3.100 3.705 -2.930 3.875 ;
        RECT -2.575 3.695 -2.405 3.865 ;
        RECT -5.840 3.390 -5.670 3.560 ;
        RECT -5.840 2.920 -5.670 3.090 ;
        RECT -5.850 2.385 -5.680 2.555 ;
        RECT -5.845 1.870 -5.675 2.040 ;
        RECT -5.845 1.130 -5.675 1.300 ;
        RECT -5.835 0.590 -5.665 0.760 ;
        RECT -5.845 -0.005 -5.675 0.165 ;
        RECT -5.845 -0.570 -5.675 -0.400 ;
        RECT -5.825 -1.230 -5.655 -1.060 ;
        RECT -5.835 -1.825 -5.665 -1.655 ;
        RECT -5.365 -1.830 -5.195 -1.660 ;
        RECT -4.840 -1.840 -4.670 -1.670 ;
        RECT -4.370 -1.845 -4.200 -1.675 ;
        RECT -3.945 -1.835 -3.775 -1.665 ;
        RECT -3.475 -1.840 -3.305 -1.670 ;
        RECT -2.950 -1.850 -2.780 -1.680 ;
        RECT 17.540 -2.360 17.710 -2.190 ;
        RECT 37.790 -2.360 37.960 -2.190 ;
        RECT 17.190 -12.205 17.360 -12.035 ;
        RECT 37.440 -12.205 37.610 -12.035 ;
        RECT 17.440 -18.960 17.610 -18.790 ;
        RECT 37.690 -18.960 37.860 -18.790 ;
      LAYER met1 ;
        RECT 15.760 14.305 17.580 15.100 ;
        RECT 8.170 14.085 17.580 14.305 ;
        RECT 8.170 6.285 8.425 14.085 ;
        RECT 15.760 13.320 17.580 14.085 ;
        RECT -2.605 6.060 8.425 6.285 ;
        RECT -2.605 3.965 -2.330 6.060 ;
        RECT 17.215 4.310 17.565 4.645 ;
        RECT 37.465 4.310 37.815 4.645 ;
        RECT -5.950 3.625 -2.330 3.965 ;
        RECT -5.950 -1.595 -5.560 3.625 ;
        RECT -5.950 -1.960 -2.355 -1.595 ;
        RECT 17.485 -3.855 17.745 -2.005 ;
        RECT 20.020 -3.855 20.380 -3.685 ;
        RECT 17.485 -4.060 20.380 -3.855 ;
        RECT 37.735 -3.855 37.995 -2.005 ;
        RECT 40.270 -3.855 40.630 -3.685 ;
        RECT 37.735 -4.060 40.630 -3.855 ;
        RECT 20.020 -9.500 40.635 -9.130 ;
        RECT 17.115 -12.290 17.465 -11.955 ;
        RECT 37.365 -12.290 37.715 -11.955 ;
        RECT 17.385 -20.455 17.645 -18.605 ;
        RECT 19.920 -20.455 20.280 -20.285 ;
        RECT 17.385 -20.660 20.280 -20.455 ;
        RECT 37.635 -20.455 37.895 -18.605 ;
        RECT 40.170 -20.455 40.530 -20.285 ;
        RECT 37.635 -20.660 40.530 -20.455 ;
      LAYER via ;
        RECT 16.030 14.380 16.290 14.640 ;
        RECT 16.555 14.405 16.815 14.665 ;
        RECT 17.075 14.405 17.335 14.665 ;
        RECT 16.030 14.060 16.290 14.320 ;
        RECT 16.555 14.085 16.815 14.345 ;
        RECT 17.075 14.085 17.335 14.345 ;
        RECT 16.030 13.740 16.290 14.000 ;
        RECT 16.555 13.765 16.815 14.025 ;
        RECT 17.075 13.765 17.335 14.025 ;
        RECT 17.265 4.335 17.525 4.595 ;
        RECT 37.525 4.350 37.785 4.610 ;
        RECT 20.065 -3.995 20.325 -3.735 ;
        RECT 40.315 -3.995 40.575 -3.735 ;
        RECT 20.065 -9.435 20.325 -9.175 ;
        RECT 40.320 -9.440 40.580 -9.180 ;
        RECT 17.140 -12.255 17.400 -11.995 ;
        RECT 37.405 -12.250 37.665 -11.990 ;
        RECT 19.965 -20.595 20.225 -20.335 ;
        RECT 40.215 -20.595 40.475 -20.335 ;
      LAYER met2 ;
        RECT 15.760 13.320 17.580 15.100 ;
        RECT 16.750 4.015 17.080 13.320 ;
        RECT 17.225 4.250 17.720 4.930 ;
        RECT 37.435 4.275 37.890 4.700 ;
        RECT 16.750 3.670 20.385 4.015 ;
        RECT 16.925 -12.500 17.500 -11.820 ;
        RECT 20.020 -20.280 20.385 3.670 ;
        RECT 40.265 -3.680 40.630 3.570 ;
        RECT 37.145 -12.700 37.885 -11.735 ;
        RECT 40.270 -20.280 40.635 -3.680 ;
        RECT 19.920 -20.660 20.385 -20.280 ;
        RECT 40.170 -20.660 40.635 -20.280 ;
      LAYER via2 ;
        RECT 16.045 14.345 16.325 14.625 ;
        RECT 16.530 14.345 16.810 14.625 ;
        RECT 17.040 14.345 17.320 14.625 ;
        RECT 16.045 13.930 16.325 14.210 ;
        RECT 16.530 13.930 16.810 14.210 ;
        RECT 17.040 13.930 17.320 14.210 ;
        RECT 16.045 13.490 16.325 13.770 ;
        RECT 16.530 13.490 16.810 13.770 ;
        RECT 17.040 13.490 17.320 13.770 ;
        RECT 17.255 4.325 17.535 4.605 ;
        RECT 37.520 4.325 37.800 4.605 ;
        RECT 16.955 -12.425 17.235 -12.145 ;
        RECT 37.395 -12.260 37.675 -11.980 ;
      LAYER met3 ;
        RECT 15.760 13.320 17.580 15.100 ;
        RECT 17.225 4.250 37.905 4.665 ;
        RECT 16.925 -12.345 17.420 -11.820 ;
        RECT 37.370 -12.345 37.700 -11.920 ;
        RECT 16.925 -12.825 37.700 -12.345 ;
        RECT 17.420 -12.830 37.700 -12.825 ;
      LAYER via3 ;
        RECT 16.025 14.325 16.345 14.645 ;
        RECT 16.510 14.325 16.830 14.645 ;
        RECT 17.020 14.325 17.340 14.645 ;
        RECT 16.025 13.910 16.345 14.230 ;
        RECT 16.510 13.910 16.830 14.230 ;
        RECT 17.020 13.910 17.340 14.230 ;
        RECT 16.025 13.470 16.345 13.790 ;
        RECT 16.510 13.470 16.830 13.790 ;
        RECT 17.020 13.470 17.340 13.790 ;
        RECT 17.235 4.305 17.555 4.625 ;
        RECT 16.935 -12.445 17.255 -12.125 ;
      LAYER met4 ;
        RECT 15.770 -14.750 17.585 165.250 ;
    END
  END vssd1
  OBS
      LAYER pwell ;
        RECT 17.120 4.170 18.130 4.790 ;
        RECT 37.370 4.170 38.380 4.790 ;
        RECT -4.860 1.875 -3.850 2.495 ;
        RECT -3.645 1.235 -2.635 2.495 ;
        RECT -2.590 -0.765 -1.580 2.495 ;
        RECT -1.555 -4.775 -0.545 2.485 ;
        RECT 14.380 -4.595 15.390 2.665 ;
        RECT 17.015 0.340 17.635 0.910 ;
        RECT 16.985 -0.160 17.665 0.340 ;
        RECT 16.985 -0.670 17.895 -0.160 ;
        RECT 16.985 -1.180 17.665 -0.670 ;
        RECT 17.015 -1.750 17.635 -1.180 ;
        RECT 18.655 -4.595 19.665 2.665 ;
        RECT 34.630 -4.595 35.640 2.665 ;
        RECT 37.265 0.340 37.885 0.910 ;
        RECT 37.235 -0.160 37.915 0.340 ;
        RECT 37.235 -0.670 38.145 -0.160 ;
        RECT 37.235 -1.180 37.915 -0.670 ;
        RECT 37.265 -1.750 37.885 -1.180 ;
        RECT 38.905 -4.595 39.915 2.665 ;
        RECT 17.020 -12.430 18.030 -11.810 ;
        RECT 37.270 -12.430 38.280 -11.810 ;
        RECT 14.280 -21.195 15.290 -13.935 ;
        RECT 16.915 -16.260 17.535 -15.690 ;
        RECT 16.885 -16.760 17.565 -16.260 ;
        RECT 16.885 -17.270 17.795 -16.760 ;
        RECT 16.885 -17.780 17.565 -17.270 ;
        RECT 16.915 -18.350 17.535 -17.780 ;
        RECT 18.555 -21.195 19.565 -13.935 ;
        RECT 34.530 -21.195 35.540 -13.935 ;
        RECT 37.165 -16.260 37.785 -15.690 ;
        RECT 37.135 -16.760 37.815 -16.260 ;
        RECT 37.135 -17.270 38.045 -16.760 ;
        RECT 37.135 -17.780 37.815 -17.270 ;
        RECT 37.165 -18.350 37.785 -17.780 ;
        RECT 38.805 -21.195 39.815 -13.935 ;
      LAYER li1 ;
        RECT 16.195 4.940 16.365 5.270 ;
        RECT 36.445 4.940 36.615 5.270 ;
        RECT -4.190 2.020 -4.020 2.350 ;
        RECT -2.975 1.400 -2.805 2.350 ;
        RECT -1.920 -0.635 -1.750 2.350 ;
        RECT -0.885 -3.000 -0.715 2.350 ;
        RECT 15.050 -2.820 15.220 2.530 ;
        RECT 15.850 1.115 16.220 4.655 ;
        RECT 17.790 4.315 17.960 4.645 ;
        RECT 17.470 1.115 17.820 3.980 ;
        RECT 16.175 0.250 17.425 0.360 ;
        RECT 16.095 0.190 17.505 0.250 ;
        RECT 16.095 -0.080 16.495 0.190 ;
        RECT 15.895 -0.590 16.145 -0.260 ;
        RECT 16.325 -0.410 16.495 -0.080 ;
        RECT 16.675 -0.060 17.005 0.020 ;
        RECT 16.675 -0.230 17.085 -0.060 ;
        RECT 17.255 -0.080 17.505 0.190 ;
        RECT 16.915 -0.250 17.085 -0.230 ;
        RECT 16.325 -0.580 16.685 -0.410 ;
        RECT 16.915 -0.420 17.345 -0.250 ;
        RECT 16.515 -0.610 16.685 -0.580 ;
        RECT 16.095 -1.030 16.345 -0.760 ;
        RECT 16.515 -0.780 17.005 -0.610 ;
        RECT 16.675 -0.860 17.005 -0.780 ;
        RECT 17.175 -0.760 17.345 -0.420 ;
        RECT 17.515 -0.580 17.765 -0.250 ;
        RECT 17.175 -1.030 17.505 -0.760 ;
        RECT 16.095 -1.090 17.505 -1.030 ;
        RECT 16.175 -1.200 17.425 -1.090 ;
        RECT 19.325 -2.820 19.495 2.530 ;
        RECT 35.300 -2.820 35.470 2.530 ;
        RECT 36.100 1.115 36.470 4.655 ;
        RECT 38.040 4.315 38.210 4.645 ;
        RECT 37.720 1.115 38.070 3.980 ;
        RECT 36.425 0.250 37.675 0.360 ;
        RECT 36.345 0.190 37.755 0.250 ;
        RECT 36.345 -0.080 36.745 0.190 ;
        RECT 36.145 -0.590 36.395 -0.260 ;
        RECT 36.575 -0.410 36.745 -0.080 ;
        RECT 36.925 -0.060 37.255 0.020 ;
        RECT 36.925 -0.230 37.335 -0.060 ;
        RECT 37.505 -0.080 37.755 0.190 ;
        RECT 37.165 -0.250 37.335 -0.230 ;
        RECT 36.575 -0.580 36.935 -0.410 ;
        RECT 37.165 -0.420 37.595 -0.250 ;
        RECT 36.765 -0.610 36.935 -0.580 ;
        RECT 36.345 -1.030 36.595 -0.760 ;
        RECT 36.765 -0.780 37.255 -0.610 ;
        RECT 36.925 -0.860 37.255 -0.780 ;
        RECT 37.425 -0.760 37.595 -0.420 ;
        RECT 37.765 -0.580 38.015 -0.250 ;
        RECT 37.425 -1.030 37.755 -0.760 ;
        RECT 36.345 -1.090 37.755 -1.030 ;
        RECT 36.425 -1.200 37.675 -1.090 ;
        RECT 39.575 -2.820 39.745 2.530 ;
        RECT 16.095 -11.660 16.265 -11.330 ;
        RECT 36.345 -11.660 36.515 -11.330 ;
        RECT 14.950 -19.420 15.120 -14.070 ;
        RECT 15.750 -15.485 16.120 -11.945 ;
        RECT 17.690 -12.285 17.860 -11.955 ;
        RECT 17.370 -15.485 17.720 -12.620 ;
        RECT 16.075 -16.350 17.325 -16.240 ;
        RECT 15.995 -16.410 17.405 -16.350 ;
        RECT 15.995 -16.680 16.395 -16.410 ;
        RECT 15.795 -17.190 16.045 -16.860 ;
        RECT 16.225 -17.010 16.395 -16.680 ;
        RECT 16.575 -16.660 16.905 -16.580 ;
        RECT 16.575 -16.830 16.985 -16.660 ;
        RECT 17.155 -16.680 17.405 -16.410 ;
        RECT 16.815 -16.850 16.985 -16.830 ;
        RECT 16.225 -17.180 16.585 -17.010 ;
        RECT 16.815 -17.020 17.245 -16.850 ;
        RECT 16.415 -17.210 16.585 -17.180 ;
        RECT 15.995 -17.630 16.245 -17.360 ;
        RECT 16.415 -17.380 16.905 -17.210 ;
        RECT 16.575 -17.460 16.905 -17.380 ;
        RECT 17.075 -17.360 17.245 -17.020 ;
        RECT 17.415 -17.180 17.665 -16.850 ;
        RECT 17.075 -17.630 17.405 -17.360 ;
        RECT 15.995 -17.690 17.405 -17.630 ;
        RECT 16.075 -17.800 17.325 -17.690 ;
        RECT 19.225 -19.420 19.395 -14.070 ;
        RECT 35.200 -19.420 35.370 -14.070 ;
        RECT 36.000 -15.485 36.370 -11.945 ;
        RECT 37.940 -12.285 38.110 -11.955 ;
        RECT 37.620 -15.485 37.970 -12.620 ;
        RECT 36.325 -16.350 37.575 -16.240 ;
        RECT 36.245 -16.410 37.655 -16.350 ;
        RECT 36.245 -16.680 36.645 -16.410 ;
        RECT 36.045 -17.190 36.295 -16.860 ;
        RECT 36.475 -17.010 36.645 -16.680 ;
        RECT 36.825 -16.660 37.155 -16.580 ;
        RECT 36.825 -16.830 37.235 -16.660 ;
        RECT 37.405 -16.680 37.655 -16.410 ;
        RECT 37.065 -16.850 37.235 -16.830 ;
        RECT 36.475 -17.180 36.835 -17.010 ;
        RECT 37.065 -17.020 37.495 -16.850 ;
        RECT 36.665 -17.210 36.835 -17.180 ;
        RECT 36.245 -17.630 36.495 -17.360 ;
        RECT 36.665 -17.380 37.155 -17.210 ;
        RECT 36.825 -17.460 37.155 -17.380 ;
        RECT 37.325 -17.360 37.495 -17.020 ;
        RECT 37.665 -17.180 37.915 -16.850 ;
        RECT 37.325 -17.630 37.655 -17.360 ;
        RECT 36.245 -17.690 37.655 -17.630 ;
        RECT 36.325 -17.800 37.575 -17.690 ;
        RECT 39.475 -19.420 39.645 -14.070 ;
      LAYER mcon ;
        RECT 16.195 5.020 16.365 5.190 ;
        RECT 36.445 5.020 36.615 5.190 ;
        RECT 15.955 4.415 16.125 4.585 ;
        RECT -4.190 2.100 -4.020 2.270 ;
        RECT -2.975 1.975 -2.805 2.145 ;
        RECT -2.975 1.615 -2.805 1.785 ;
        RECT -1.920 1.800 -1.750 1.970 ;
        RECT -1.920 1.440 -1.750 1.610 ;
        RECT -1.920 1.080 -1.750 1.250 ;
        RECT -1.920 0.720 -1.750 0.890 ;
        RECT -1.920 0.360 -1.750 0.530 ;
        RECT -1.920 0.000 -1.750 0.170 ;
        RECT -1.920 -0.360 -1.750 -0.190 ;
        RECT -0.885 1.960 -0.715 2.130 ;
        RECT -0.885 1.600 -0.715 1.770 ;
        RECT -0.885 1.240 -0.715 1.410 ;
        RECT -0.885 0.880 -0.715 1.050 ;
        RECT -0.885 0.520 -0.715 0.690 ;
        RECT -0.885 0.160 -0.715 0.330 ;
        RECT -0.885 -0.200 -0.715 -0.030 ;
        RECT -0.885 -0.560 -0.715 -0.390 ;
        RECT -0.885 -0.920 -0.715 -0.750 ;
        RECT -0.885 -1.280 -0.715 -1.110 ;
        RECT -0.885 -1.640 -0.715 -1.470 ;
        RECT -0.885 -2.000 -0.715 -1.830 ;
        RECT -0.885 -2.360 -0.715 -2.190 ;
        RECT -0.885 -2.720 -0.715 -2.550 ;
        RECT 15.050 2.140 15.220 2.310 ;
        RECT 15.050 1.780 15.220 1.950 ;
        RECT 15.050 1.420 15.220 1.590 ;
        RECT 15.050 1.060 15.220 1.230 ;
        RECT 17.790 4.395 17.960 4.565 ;
        RECT 36.205 4.395 36.375 4.565 ;
        RECT 15.950 1.225 16.120 1.395 ;
        RECT 17.550 3.760 17.720 3.930 ;
        RECT 17.535 1.220 17.705 1.390 ;
        RECT 19.325 2.140 19.495 2.310 ;
        RECT 19.325 1.780 19.495 1.950 ;
        RECT 19.325 1.420 19.495 1.590 ;
        RECT 15.050 0.700 15.220 0.870 ;
        RECT 15.050 0.340 15.220 0.510 ;
        RECT 19.325 1.060 19.495 1.230 ;
        RECT 19.325 0.700 19.495 0.870 ;
        RECT 19.325 0.340 19.495 0.510 ;
        RECT 15.050 -0.020 15.220 0.150 ;
        RECT 15.050 -0.380 15.220 -0.210 ;
        RECT 15.050 -0.740 15.220 -0.570 ;
        RECT 15.975 -0.510 16.145 -0.340 ;
        RECT 19.325 -0.020 19.495 0.150 ;
        RECT 15.050 -1.100 15.220 -0.930 ;
        RECT 17.515 -0.500 17.685 -0.330 ;
        RECT 19.325 -0.380 19.495 -0.210 ;
        RECT 19.325 -0.740 19.495 -0.570 ;
        RECT 19.325 -1.100 19.495 -0.930 ;
        RECT 15.050 -1.460 15.220 -1.290 ;
        RECT 15.050 -1.820 15.220 -1.650 ;
        RECT 15.050 -2.180 15.220 -2.010 ;
        RECT 15.050 -2.540 15.220 -2.370 ;
        RECT 19.325 -1.460 19.495 -1.290 ;
        RECT 19.325 -1.820 19.495 -1.650 ;
        RECT 19.325 -2.180 19.495 -2.010 ;
        RECT 19.325 -2.540 19.495 -2.370 ;
        RECT 35.300 2.140 35.470 2.310 ;
        RECT 35.300 1.780 35.470 1.950 ;
        RECT 35.300 1.420 35.470 1.590 ;
        RECT 35.300 1.060 35.470 1.230 ;
        RECT 38.040 4.395 38.210 4.565 ;
        RECT 36.200 1.225 36.370 1.395 ;
        RECT 37.800 3.755 37.970 3.925 ;
        RECT 37.785 1.220 37.955 1.390 ;
        RECT 39.575 2.140 39.745 2.310 ;
        RECT 39.575 1.780 39.745 1.950 ;
        RECT 39.575 1.420 39.745 1.590 ;
        RECT 35.300 0.700 35.470 0.870 ;
        RECT 35.300 0.340 35.470 0.510 ;
        RECT 39.575 1.060 39.745 1.230 ;
        RECT 39.575 0.700 39.745 0.870 ;
        RECT 39.575 0.340 39.745 0.510 ;
        RECT 35.300 -0.020 35.470 0.150 ;
        RECT 35.300 -0.380 35.470 -0.210 ;
        RECT 35.300 -0.740 35.470 -0.570 ;
        RECT 36.225 -0.510 36.395 -0.340 ;
        RECT 39.575 -0.020 39.745 0.150 ;
        RECT 35.300 -1.100 35.470 -0.930 ;
        RECT 37.765 -0.500 37.935 -0.330 ;
        RECT 39.575 -0.380 39.745 -0.210 ;
        RECT 39.575 -0.740 39.745 -0.570 ;
        RECT 39.575 -1.100 39.745 -0.930 ;
        RECT 35.300 -1.460 35.470 -1.290 ;
        RECT 35.300 -1.820 35.470 -1.650 ;
        RECT 35.300 -2.180 35.470 -2.010 ;
        RECT 35.300 -2.540 35.470 -2.370 ;
        RECT 39.575 -1.460 39.745 -1.290 ;
        RECT 39.575 -1.820 39.745 -1.650 ;
        RECT 39.575 -2.180 39.745 -2.010 ;
        RECT 39.575 -2.540 39.745 -2.370 ;
        RECT 16.095 -11.580 16.265 -11.410 ;
        RECT 36.345 -11.580 36.515 -11.410 ;
        RECT 15.855 -12.185 16.025 -12.015 ;
        RECT 14.950 -14.460 15.120 -14.290 ;
        RECT 14.950 -14.820 15.120 -14.650 ;
        RECT 14.950 -15.180 15.120 -15.010 ;
        RECT 14.950 -15.540 15.120 -15.370 ;
        RECT 17.690 -12.205 17.860 -12.035 ;
        RECT 36.105 -12.190 36.275 -12.020 ;
        RECT 15.850 -15.375 16.020 -15.205 ;
        RECT 17.450 -12.840 17.620 -12.670 ;
        RECT 17.435 -15.380 17.605 -15.210 ;
        RECT 19.225 -14.460 19.395 -14.290 ;
        RECT 19.225 -14.820 19.395 -14.650 ;
        RECT 19.225 -15.180 19.395 -15.010 ;
        RECT 14.950 -15.900 15.120 -15.730 ;
        RECT 14.950 -16.260 15.120 -16.090 ;
        RECT 19.225 -15.540 19.395 -15.370 ;
        RECT 19.225 -15.900 19.395 -15.730 ;
        RECT 19.225 -16.260 19.395 -16.090 ;
        RECT 14.950 -16.620 15.120 -16.450 ;
        RECT 14.950 -16.980 15.120 -16.810 ;
        RECT 14.950 -17.340 15.120 -17.170 ;
        RECT 15.875 -17.110 16.045 -16.940 ;
        RECT 19.225 -16.620 19.395 -16.450 ;
        RECT 14.950 -17.700 15.120 -17.530 ;
        RECT 17.415 -17.100 17.585 -16.930 ;
        RECT 19.225 -16.980 19.395 -16.810 ;
        RECT 19.225 -17.340 19.395 -17.170 ;
        RECT 19.225 -17.700 19.395 -17.530 ;
        RECT 14.950 -18.060 15.120 -17.890 ;
        RECT 14.950 -18.420 15.120 -18.250 ;
        RECT 14.950 -18.780 15.120 -18.610 ;
        RECT 14.950 -19.140 15.120 -18.970 ;
        RECT 19.225 -18.060 19.395 -17.890 ;
        RECT 19.225 -18.420 19.395 -18.250 ;
        RECT 19.225 -18.780 19.395 -18.610 ;
        RECT 19.225 -19.140 19.395 -18.970 ;
        RECT 35.200 -14.460 35.370 -14.290 ;
        RECT 35.200 -14.820 35.370 -14.650 ;
        RECT 35.200 -15.180 35.370 -15.010 ;
        RECT 35.200 -15.540 35.370 -15.370 ;
        RECT 37.940 -12.205 38.110 -12.035 ;
        RECT 36.100 -15.375 36.270 -15.205 ;
        RECT 37.700 -12.840 37.870 -12.670 ;
        RECT 37.685 -15.380 37.855 -15.210 ;
        RECT 39.475 -14.460 39.645 -14.290 ;
        RECT 39.475 -14.820 39.645 -14.650 ;
        RECT 39.475 -15.180 39.645 -15.010 ;
        RECT 35.200 -15.900 35.370 -15.730 ;
        RECT 35.200 -16.260 35.370 -16.090 ;
        RECT 39.475 -15.540 39.645 -15.370 ;
        RECT 39.475 -15.900 39.645 -15.730 ;
        RECT 39.475 -16.260 39.645 -16.090 ;
        RECT 35.200 -16.620 35.370 -16.450 ;
        RECT 35.200 -16.980 35.370 -16.810 ;
        RECT 35.200 -17.340 35.370 -17.170 ;
        RECT 36.125 -17.110 36.295 -16.940 ;
        RECT 39.475 -16.620 39.645 -16.450 ;
        RECT 35.200 -17.700 35.370 -17.530 ;
        RECT 37.665 -17.100 37.835 -16.930 ;
        RECT 39.475 -16.980 39.645 -16.810 ;
        RECT 39.475 -17.340 39.645 -17.170 ;
        RECT 39.475 -17.700 39.645 -17.530 ;
        RECT 35.200 -18.060 35.370 -17.890 ;
        RECT 35.200 -18.420 35.370 -18.250 ;
        RECT 35.200 -18.780 35.370 -18.610 ;
        RECT 35.200 -19.140 35.370 -18.970 ;
        RECT 39.475 -18.060 39.645 -17.890 ;
        RECT 39.475 -18.420 39.645 -18.250 ;
        RECT 39.475 -18.780 39.645 -18.610 ;
        RECT 39.475 -19.140 39.645 -18.970 ;
      LAYER met1 ;
        RECT 16.165 4.960 16.395 5.270 ;
        RECT 36.415 4.960 36.645 5.270 ;
        RECT 16.210 4.795 16.350 4.960 ;
        RECT 36.460 4.795 36.600 4.960 ;
        RECT 15.955 4.655 16.350 4.795 ;
        RECT 36.205 4.655 36.600 4.795 ;
        RECT 15.850 4.265 16.220 4.655 ;
        RECT 17.760 4.335 17.990 4.645 ;
        RECT 17.805 4.170 17.945 4.335 ;
        RECT 36.100 4.275 36.470 4.655 ;
        RECT 38.010 4.335 38.240 4.645 ;
        RECT 38.055 4.170 38.195 4.335 ;
        RECT 17.550 4.030 17.945 4.170 ;
        RECT 37.800 4.030 38.195 4.170 ;
        RECT 17.470 3.670 17.820 4.030 ;
        RECT 37.720 3.670 38.070 4.030 ;
        RECT -4.530 2.950 -4.210 3.210 ;
        RECT -3.315 2.950 -2.995 3.210 ;
        RECT -2.260 2.950 -1.940 3.210 ;
        RECT -1.225 2.950 -0.905 3.210 ;
        RECT 14.710 3.130 15.030 3.390 ;
        RECT 18.985 3.130 19.305 3.390 ;
        RECT 34.960 3.130 35.280 3.390 ;
        RECT 39.235 3.130 39.555 3.390 ;
        RECT -4.430 2.635 -4.270 2.950 ;
        RECT -3.215 2.635 -3.055 2.950 ;
        RECT -2.160 2.635 -2.000 2.950 ;
        RECT -1.125 2.635 -0.965 2.950 ;
        RECT 14.810 2.815 14.970 3.130 ;
        RECT 19.085 2.815 19.245 3.130 ;
        RECT 35.060 2.815 35.220 3.130 ;
        RECT 39.335 2.815 39.495 3.130 ;
        RECT 14.810 2.675 15.205 2.815 ;
        RECT 19.085 2.675 19.480 2.815 ;
        RECT 35.060 2.675 35.455 2.815 ;
        RECT 39.335 2.675 39.730 2.815 ;
        RECT -4.430 2.495 -4.035 2.635 ;
        RECT -3.215 2.495 -2.820 2.635 ;
        RECT -2.160 2.495 -1.765 2.635 ;
        RECT -1.125 2.495 -0.730 2.635 ;
        RECT 15.065 2.510 15.205 2.675 ;
        RECT 19.340 2.510 19.480 2.675 ;
        RECT 35.315 2.510 35.455 2.675 ;
        RECT 39.590 2.510 39.730 2.675 ;
        RECT -4.175 2.330 -4.035 2.495 ;
        RECT -2.960 2.330 -2.820 2.495 ;
        RECT -1.905 2.330 -1.765 2.495 ;
        RECT -0.870 2.330 -0.730 2.495 ;
        RECT -4.220 2.020 -3.990 2.330 ;
        RECT -3.005 1.395 -2.775 2.330 ;
        RECT -1.950 -0.635 -1.720 2.330 ;
        RECT -0.915 -3.000 -0.685 2.330 ;
        RECT 15.020 -2.820 15.250 2.510 ;
        RECT 15.915 0.360 16.175 1.490 ;
        RECT 17.505 0.780 17.745 1.490 ;
        RECT 15.915 0.040 16.235 0.360 ;
        RECT 15.915 -0.280 16.175 0.040 ;
        RECT 17.485 -0.260 17.745 0.780 ;
        RECT 15.915 -0.570 16.205 -0.280 ;
        RECT 15.915 -1.620 16.175 -0.570 ;
        RECT 17.425 -0.580 17.745 -0.260 ;
        RECT 17.485 -1.620 17.745 -0.580 ;
        RECT 19.295 -2.820 19.525 2.510 ;
        RECT 35.270 -2.820 35.500 2.510 ;
        RECT 36.165 0.360 36.425 1.490 ;
        RECT 37.755 0.780 37.995 1.490 ;
        RECT 36.165 0.040 36.485 0.360 ;
        RECT 36.165 -0.280 36.425 0.040 ;
        RECT 37.735 -0.260 37.995 0.780 ;
        RECT 36.165 -0.570 36.455 -0.280 ;
        RECT 36.165 -1.620 36.425 -0.570 ;
        RECT 37.675 -0.580 37.995 -0.260 ;
        RECT 37.735 -1.620 37.995 -0.580 ;
        RECT 39.545 -2.820 39.775 2.510 ;
        RECT 16.065 -11.640 16.295 -11.330 ;
        RECT 36.315 -11.640 36.545 -11.330 ;
        RECT 16.110 -11.805 16.250 -11.640 ;
        RECT 36.360 -11.805 36.500 -11.640 ;
        RECT 15.855 -11.945 16.250 -11.805 ;
        RECT 36.105 -11.945 36.500 -11.805 ;
        RECT 15.750 -12.295 16.120 -11.945 ;
        RECT 17.660 -12.265 17.890 -11.955 ;
        RECT 17.705 -12.430 17.845 -12.265 ;
        RECT 36.000 -12.275 36.370 -11.945 ;
        RECT 37.910 -12.265 38.140 -11.955 ;
        RECT 37.955 -12.430 38.095 -12.265 ;
        RECT 17.450 -12.570 17.845 -12.430 ;
        RECT 37.700 -12.570 38.095 -12.430 ;
        RECT 17.370 -12.985 17.720 -12.570 ;
        RECT 37.620 -12.920 37.970 -12.570 ;
        RECT 14.610 -13.470 14.930 -13.210 ;
        RECT 18.885 -13.470 19.205 -13.210 ;
        RECT 34.860 -13.470 35.180 -13.210 ;
        RECT 39.135 -13.470 39.455 -13.210 ;
        RECT 14.710 -13.785 14.870 -13.470 ;
        RECT 18.985 -13.785 19.145 -13.470 ;
        RECT 34.960 -13.785 35.120 -13.470 ;
        RECT 39.235 -13.785 39.395 -13.470 ;
        RECT 14.710 -13.925 15.105 -13.785 ;
        RECT 18.985 -13.925 19.380 -13.785 ;
        RECT 34.960 -13.925 35.355 -13.785 ;
        RECT 39.235 -13.925 39.630 -13.785 ;
        RECT 14.965 -14.090 15.105 -13.925 ;
        RECT 19.240 -14.090 19.380 -13.925 ;
        RECT 35.215 -14.090 35.355 -13.925 ;
        RECT 39.490 -14.090 39.630 -13.925 ;
        RECT 14.920 -19.420 15.150 -14.090 ;
        RECT 15.815 -16.240 16.075 -15.110 ;
        RECT 17.405 -15.820 17.645 -15.110 ;
        RECT 15.815 -16.560 16.135 -16.240 ;
        RECT 15.815 -16.880 16.075 -16.560 ;
        RECT 17.385 -16.860 17.645 -15.820 ;
        RECT 15.815 -17.170 16.105 -16.880 ;
        RECT 15.815 -18.220 16.075 -17.170 ;
        RECT 17.325 -17.180 17.645 -16.860 ;
        RECT 17.385 -18.220 17.645 -17.180 ;
        RECT 19.195 -19.420 19.425 -14.090 ;
        RECT 35.170 -19.420 35.400 -14.090 ;
        RECT 36.065 -16.240 36.325 -15.110 ;
        RECT 37.655 -15.820 37.895 -15.110 ;
        RECT 36.065 -16.560 36.385 -16.240 ;
        RECT 36.065 -16.880 36.325 -16.560 ;
        RECT 37.635 -16.860 37.895 -15.820 ;
        RECT 36.065 -17.170 36.355 -16.880 ;
        RECT 36.065 -18.220 36.325 -17.170 ;
        RECT 37.575 -17.180 37.895 -16.860 ;
        RECT 37.635 -18.220 37.895 -17.180 ;
        RECT 39.445 -19.420 39.675 -14.090 ;
      LAYER via ;
        RECT 15.945 0.070 16.205 0.330 ;
        RECT 17.455 -0.550 17.715 -0.290 ;
        RECT 36.195 0.070 36.455 0.330 ;
        RECT 37.705 -0.550 37.965 -0.290 ;
        RECT 15.845 -16.530 16.105 -16.270 ;
        RECT 17.355 -17.150 17.615 -16.890 ;
        RECT 36.095 -16.530 36.355 -16.270 ;
        RECT 37.605 -17.150 37.865 -16.890 ;
      LAYER met2 ;
        RECT 15.895 0.040 17.765 0.360 ;
        RECT 36.145 0.040 38.015 0.360 ;
        RECT 15.895 -0.580 17.765 -0.260 ;
        RECT 36.145 -0.580 38.015 -0.260 ;
        RECT 15.895 -1.200 17.765 -0.880 ;
        RECT 36.145 -1.200 38.015 -0.880 ;
        RECT 15.795 -16.560 17.665 -16.240 ;
        RECT 36.045 -16.560 37.915 -16.240 ;
        RECT 15.795 -17.180 17.665 -16.860 ;
        RECT 36.045 -17.180 37.915 -16.860 ;
        RECT 15.795 -17.800 17.665 -17.480 ;
        RECT 36.045 -17.800 37.915 -17.480 ;
  END
END rram_test
END LIBRARY


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO 1T1R_700U
  CLASS BLOCK ;
  FOREIGN 1T1R_700U ;
  ORIGIN 0.920 13.910 ;
  SIZE 1.010 BY 8.375 ;
  PIN G
    ANTENNAGATEAREA 1.050000 ;
    PORT
      LAYER li1 ;
        RECT -0.570 -13.910 -0.215 -13.625 ;
    END
  END G
  PIN S
    ANTENNADIFFAREA 2.100000 ;
    PORT
      LAYER li1 ;
        RECT -0.750 -11.805 -0.580 -6.455 ;
      LAYER mcon ;
        RECT -0.750 -6.840 -0.580 -6.670 ;
        RECT -0.750 -7.200 -0.580 -7.030 ;
        RECT -0.750 -7.560 -0.580 -7.390 ;
        RECT -0.750 -7.920 -0.580 -7.750 ;
        RECT -0.750 -8.280 -0.580 -8.110 ;
        RECT -0.750 -8.640 -0.580 -8.470 ;
        RECT -0.750 -9.000 -0.580 -8.830 ;
        RECT -0.750 -9.360 -0.580 -9.190 ;
        RECT -0.750 -9.720 -0.580 -9.550 ;
        RECT -0.750 -10.080 -0.580 -9.910 ;
        RECT -0.750 -10.440 -0.580 -10.270 ;
        RECT -0.750 -10.800 -0.580 -10.630 ;
        RECT -0.750 -11.160 -0.580 -10.990 ;
        RECT -0.750 -11.520 -0.580 -11.350 ;
      LAYER met1 ;
        RECT -0.795 -11.805 -0.475 -6.450 ;
      LAYER via ;
        RECT -0.765 -6.915 -0.505 -6.655 ;
        RECT -0.765 -7.235 -0.505 -6.975 ;
        RECT -0.765 -7.555 -0.505 -7.295 ;
        RECT -0.765 -7.875 -0.505 -7.615 ;
        RECT -0.765 -8.195 -0.505 -7.935 ;
        RECT -0.765 -8.515 -0.505 -8.255 ;
        RECT -0.765 -8.835 -0.505 -8.575 ;
        RECT -0.765 -9.155 -0.505 -8.895 ;
        RECT -0.765 -9.475 -0.505 -9.215 ;
        RECT -0.765 -9.795 -0.505 -9.535 ;
        RECT -0.765 -10.115 -0.505 -9.855 ;
        RECT -0.765 -10.435 -0.505 -10.175 ;
        RECT -0.765 -10.755 -0.505 -10.495 ;
        RECT -0.765 -11.075 -0.505 -10.815 ;
        RECT -0.765 -11.395 -0.505 -11.135 ;
        RECT -0.765 -11.715 -0.505 -11.455 ;
      LAYER met2 ;
        RECT -0.795 -11.800 -0.475 -6.450 ;
    END
  END S
  OBS
      LAYER pwell ;
        RECT -0.920 -13.580 0.090 -6.320 ;
      LAYER li1 ;
        RECT -0.250 -11.805 -0.080 -6.455 ;
      LAYER mcon ;
        RECT -0.250 -6.845 -0.080 -6.675 ;
        RECT -0.250 -7.205 -0.080 -7.035 ;
        RECT -0.250 -7.565 -0.080 -7.395 ;
        RECT -0.250 -7.925 -0.080 -7.755 ;
        RECT -0.250 -8.285 -0.080 -8.115 ;
        RECT -0.250 -8.645 -0.080 -8.475 ;
        RECT -0.250 -9.005 -0.080 -8.835 ;
        RECT -0.250 -9.365 -0.080 -9.195 ;
        RECT -0.250 -9.725 -0.080 -9.555 ;
        RECT -0.250 -10.085 -0.080 -9.915 ;
        RECT -0.250 -10.445 -0.080 -10.275 ;
        RECT -0.250 -10.805 -0.080 -10.635 ;
        RECT -0.250 -11.165 -0.080 -10.995 ;
        RECT -0.250 -11.525 -0.080 -11.355 ;
      LAYER met1 ;
        RECT -0.590 -5.855 -0.270 -5.595 ;
        RECT -0.490 -6.170 -0.330 -5.855 ;
        RECT -0.490 -6.310 -0.095 -6.170 ;
        RECT -0.235 -6.475 -0.095 -6.310 ;
        RECT -0.280 -11.805 -0.050 -6.475 ;
  END
END 1T1R_700U
MACRO array
  CLASS BLOCK ;
  FOREIGN array ;
  ORIGIN 6.960 16.895 ;
  SIZE 34.920 BY 29.775 ;
  PIN re_wl1
    ANTENNAGATEAREA 4.200000 ;
    PORT
      LAYER li1 ;
        RECT -6.960 -16.035 5.110 -15.865 ;
        RECT 13.290 -16.035 22.200 -15.865 ;
        RECT -3.080 -16.715 -2.725 -16.035 ;
        RECT 1.195 -16.715 1.550 -16.035 ;
        RECT 17.170 -16.715 17.525 -16.035 ;
        RECT 21.445 -16.715 21.800 -16.035 ;
      LAYER mcon ;
        RECT 4.855 -16.035 5.025 -15.865 ;
        RECT 13.400 -16.035 13.570 -15.865 ;
      LAYER met1 ;
        RECT 4.745 -16.185 13.655 -15.820 ;
    END
  END re_wl1
  PIN wl1
    ANTENNAGATEAREA 0.216000 ;
    PORT
      LAYER li1 ;
        RECT -2.420 -15.405 -2.105 -14.850 ;
        RECT 17.830 -15.405 18.145 -14.850 ;
        RECT -6.960 -15.575 5.110 -15.405 ;
        RECT 13.290 -15.575 22.200 -15.405 ;
      LAYER mcon ;
        RECT 4.855 -15.575 5.025 -15.405 ;
        RECT 13.400 -15.575 13.570 -15.405 ;
      LAYER met1 ;
        RECT 4.745 -15.620 13.655 -15.230 ;
    END
  END wl1
  PIN wl0
    ANTENNAGATEAREA 0.216000 ;
    PORT
      LAYER li1 ;
        RECT -2.320 1.195 -2.005 1.750 ;
        RECT 17.930 1.195 18.245 1.750 ;
        RECT -6.860 1.025 5.015 1.195 ;
        RECT 13.390 1.025 22.200 1.195 ;
      LAYER mcon ;
        RECT 4.760 1.025 4.930 1.195 ;
        RECT 13.500 1.025 13.670 1.195 ;
      LAYER met1 ;
        RECT 4.650 0.980 13.755 1.370 ;
    END
  END wl0
  PIN re_wl0
    ANTENNAGATEAREA 4.200000 ;
    PORT
      LAYER li1 ;
        RECT -6.860 0.565 5.015 0.735 ;
        RECT 13.390 0.565 22.200 0.735 ;
        RECT -2.980 -0.115 -2.625 0.565 ;
        RECT 1.295 -0.115 1.650 0.565 ;
        RECT 17.270 -0.115 17.625 0.565 ;
        RECT 21.545 -0.115 21.900 0.565 ;
      LAYER mcon ;
        RECT 4.760 0.565 4.930 0.735 ;
        RECT 13.500 0.565 13.670 0.735 ;
      LAYER met1 ;
        RECT 4.650 0.415 13.755 0.780 ;
    END
  END re_wl0
  PIN re_br1
    ANTENNADIFFAREA 4.200000 ;
    PORT
      LAYER li1 ;
        RECT 21.365 1.990 21.535 7.340 ;
        RECT 21.265 -14.610 21.435 -9.260 ;
      LAYER mcon ;
        RECT 21.365 6.955 21.535 7.125 ;
        RECT 21.365 6.595 21.535 6.765 ;
        RECT 21.365 6.235 21.535 6.405 ;
        RECT 21.365 5.875 21.535 6.045 ;
        RECT 21.365 5.515 21.535 5.685 ;
        RECT 21.365 5.155 21.535 5.325 ;
        RECT 21.365 4.795 21.535 4.965 ;
        RECT 21.365 4.435 21.535 4.605 ;
        RECT 21.365 4.075 21.535 4.245 ;
        RECT 21.365 3.715 21.535 3.885 ;
        RECT 21.365 3.355 21.535 3.525 ;
        RECT 21.365 2.995 21.535 3.165 ;
        RECT 21.365 2.635 21.535 2.805 ;
        RECT 21.365 2.275 21.535 2.445 ;
        RECT 21.265 -9.645 21.435 -9.475 ;
        RECT 21.265 -10.005 21.435 -9.835 ;
        RECT 21.265 -10.365 21.435 -10.195 ;
        RECT 21.265 -10.725 21.435 -10.555 ;
        RECT 21.265 -11.085 21.435 -10.915 ;
        RECT 21.265 -11.445 21.435 -11.275 ;
        RECT 21.265 -11.805 21.435 -11.635 ;
        RECT 21.265 -12.165 21.435 -11.995 ;
        RECT 21.265 -12.525 21.435 -12.355 ;
        RECT 21.265 -12.885 21.435 -12.715 ;
        RECT 21.265 -13.245 21.435 -13.075 ;
        RECT 21.265 -13.605 21.435 -13.435 ;
        RECT 21.265 -13.965 21.435 -13.795 ;
        RECT 21.265 -14.325 21.435 -14.155 ;
      LAYER met1 ;
        RECT 21.320 1.730 21.640 7.345 ;
        RECT 21.320 1.525 24.235 1.730 ;
        RECT 23.955 -0.160 24.235 1.525 ;
        RECT 21.220 -14.870 21.540 -9.255 ;
        RECT 21.220 -15.075 24.135 -14.870 ;
        RECT 23.855 -16.760 24.135 -15.075 ;
      LAYER via ;
        RECT 21.350 6.880 21.610 7.140 ;
        RECT 21.350 6.560 21.610 6.820 ;
        RECT 21.350 6.240 21.610 6.500 ;
        RECT 21.350 5.920 21.610 6.180 ;
        RECT 21.350 5.600 21.610 5.860 ;
        RECT 21.350 5.280 21.610 5.540 ;
        RECT 21.350 4.960 21.610 5.220 ;
        RECT 21.350 4.640 21.610 4.900 ;
        RECT 21.350 4.320 21.610 4.580 ;
        RECT 21.350 4.000 21.610 4.260 ;
        RECT 21.350 3.680 21.610 3.940 ;
        RECT 21.350 3.360 21.610 3.620 ;
        RECT 21.350 3.040 21.610 3.300 ;
        RECT 21.350 2.720 21.610 2.980 ;
        RECT 21.350 2.400 21.610 2.660 ;
        RECT 21.350 2.080 21.610 2.340 ;
        RECT 23.960 -0.100 24.220 0.160 ;
        RECT 21.250 -9.720 21.510 -9.460 ;
        RECT 21.250 -10.040 21.510 -9.780 ;
        RECT 21.250 -10.360 21.510 -10.100 ;
        RECT 21.250 -10.680 21.510 -10.420 ;
        RECT 21.250 -11.000 21.510 -10.740 ;
        RECT 21.250 -11.320 21.510 -11.060 ;
        RECT 21.250 -11.640 21.510 -11.380 ;
        RECT 21.250 -11.960 21.510 -11.700 ;
        RECT 21.250 -12.280 21.510 -12.020 ;
        RECT 21.250 -12.600 21.510 -12.340 ;
        RECT 21.250 -12.920 21.510 -12.660 ;
        RECT 21.250 -13.240 21.510 -12.980 ;
        RECT 21.250 -13.560 21.510 -13.300 ;
        RECT 21.250 -13.880 21.510 -13.620 ;
        RECT 21.250 -14.200 21.510 -13.940 ;
        RECT 21.250 -14.520 21.510 -14.260 ;
        RECT 23.860 -16.700 24.120 -16.440 ;
      LAYER met2 ;
        RECT 21.320 1.995 21.640 7.345 ;
        RECT 21.220 -14.605 21.540 -9.255 ;
        RECT 23.730 -16.370 24.235 0.230 ;
        RECT 23.630 -16.760 24.235 -16.370 ;
    END
  END re_br1
  PIN br1
    ANTENNADIFFAREA 0.244800 ;
    PORT
      LAYER li1 ;
        RECT 18.705 3.190 20.045 3.440 ;
        RECT 18.605 -13.410 19.945 -13.160 ;
      LAYER mcon ;
        RECT 19.555 3.230 19.725 3.400 ;
        RECT 19.455 -13.370 19.625 -13.200 ;
      LAYER met1 ;
        RECT 19.495 7.650 20.385 8.230 ;
        RECT 19.495 5.590 19.785 7.650 ;
        RECT 19.505 3.460 19.765 5.590 ;
        RECT 19.495 3.190 19.785 3.460 ;
        RECT 19.505 0.610 19.765 3.190 ;
        RECT 23.200 0.610 23.475 0.830 ;
        RECT 19.505 0.405 23.475 0.610 ;
        RECT 19.505 0.400 19.765 0.405 ;
        RECT 19.395 -8.950 20.285 -8.370 ;
        RECT 19.395 -11.010 19.685 -8.950 ;
        RECT 19.405 -13.140 19.665 -11.010 ;
        RECT 19.395 -13.410 19.685 -13.140 ;
        RECT 19.405 -15.990 19.665 -13.410 ;
        RECT 23.100 -15.990 23.375 -15.770 ;
        RECT 19.405 -16.195 23.375 -15.990 ;
        RECT 19.405 -16.200 19.665 -16.195 ;
      LAYER via ;
        RECT 19.965 7.800 20.225 8.060 ;
        RECT 23.205 0.460 23.465 0.720 ;
        RECT 19.865 -8.800 20.125 -8.540 ;
        RECT 23.105 -16.140 23.365 -15.880 ;
      LAYER met2 ;
        RECT 19.790 7.960 21.525 8.230 ;
        RECT 19.790 7.655 20.380 7.960 ;
        RECT 19.690 -8.640 21.425 -8.370 ;
        RECT 19.690 -8.945 20.280 -8.640 ;
        RECT 23.195 -15.765 23.485 0.835 ;
        RECT 23.095 -16.190 23.485 -15.765 ;
    END
  END br1
  PIN gnd
    PORT
      LAYER li1 ;
        RECT 20.030 2.305 20.290 2.885 ;
        RECT 19.930 -14.295 20.190 -13.715 ;
      LAYER mcon ;
        RECT 20.080 2.450 20.250 2.620 ;
        RECT 19.980 -14.150 20.150 -13.980 ;
      LAYER met1 ;
        RECT 20.025 0.955 20.285 2.805 ;
        RECT 22.560 0.955 22.920 1.125 ;
        RECT 20.025 0.750 22.920 0.955 ;
        RECT 19.925 -15.645 20.185 -13.795 ;
        RECT 22.460 -15.645 22.820 -15.475 ;
        RECT 19.925 -15.850 22.820 -15.645 ;
      LAYER via ;
        RECT 22.605 0.815 22.865 1.075 ;
        RECT 22.505 -15.785 22.765 -15.525 ;
      LAYER met2 ;
        RECT 22.560 -15.470 22.925 1.130 ;
        RECT 22.460 -15.850 22.925 -15.470 ;
    END
    PORT
      LAYER li1 ;
        RECT -0.220 2.305 0.040 2.885 ;
        RECT -0.320 -14.295 -0.060 -13.715 ;
      LAYER mcon ;
        RECT -0.170 2.450 0.000 2.620 ;
        RECT -0.270 -14.150 -0.100 -13.980 ;
      LAYER met1 ;
        RECT -0.225 0.955 0.035 2.805 ;
        RECT 2.310 0.955 2.670 1.125 ;
        RECT -0.225 0.750 2.670 0.955 ;
        RECT -0.325 -15.645 -0.065 -13.795 ;
        RECT 2.210 -15.645 2.570 -15.475 ;
        RECT -0.325 -15.850 2.570 -15.645 ;
      LAYER via ;
        RECT 2.355 0.815 2.615 1.075 ;
        RECT 2.255 -15.785 2.515 -15.525 ;
      LAYER met2 ;
        RECT 2.310 -15.470 2.675 1.130 ;
        RECT 2.210 -15.850 2.675 -15.470 ;
    END
  END gnd
  PIN re_bl1
    ANTENNADIFFAREA 4.200000 ;
    PORT
      LAYER li1 ;
        RECT 17.090 1.990 17.260 7.340 ;
        RECT 16.990 -14.610 17.160 -9.260 ;
      LAYER mcon ;
        RECT 17.090 6.955 17.260 7.125 ;
        RECT 17.090 6.595 17.260 6.765 ;
        RECT 17.090 6.235 17.260 6.405 ;
        RECT 17.090 5.875 17.260 6.045 ;
        RECT 17.090 5.515 17.260 5.685 ;
        RECT 17.090 5.155 17.260 5.325 ;
        RECT 17.090 4.795 17.260 4.965 ;
        RECT 17.090 4.435 17.260 4.605 ;
        RECT 17.090 4.075 17.260 4.245 ;
        RECT 17.090 3.715 17.260 3.885 ;
        RECT 17.090 3.355 17.260 3.525 ;
        RECT 17.090 2.995 17.260 3.165 ;
        RECT 17.090 2.635 17.260 2.805 ;
        RECT 17.090 2.275 17.260 2.445 ;
        RECT 16.990 -9.645 17.160 -9.475 ;
        RECT 16.990 -10.005 17.160 -9.835 ;
        RECT 16.990 -10.365 17.160 -10.195 ;
        RECT 16.990 -10.725 17.160 -10.555 ;
        RECT 16.990 -11.085 17.160 -10.915 ;
        RECT 16.990 -11.445 17.160 -11.275 ;
        RECT 16.990 -11.805 17.160 -11.635 ;
        RECT 16.990 -12.165 17.160 -11.995 ;
        RECT 16.990 -12.525 17.160 -12.355 ;
        RECT 16.990 -12.885 17.160 -12.715 ;
        RECT 16.990 -13.245 17.160 -13.075 ;
        RECT 16.990 -13.605 17.160 -13.435 ;
        RECT 16.990 -13.965 17.160 -13.795 ;
        RECT 16.990 -14.325 17.160 -14.155 ;
      LAYER met1 ;
        RECT 17.045 2.345 17.365 7.345 ;
        RECT 14.785 2.030 17.365 2.345 ;
        RECT 14.785 -0.115 15.150 2.030 ;
        RECT 17.045 1.990 17.365 2.030 ;
        RECT 16.945 -14.255 17.265 -9.255 ;
        RECT 14.685 -14.570 17.265 -14.255 ;
        RECT 14.685 -16.715 15.050 -14.570 ;
        RECT 16.945 -14.610 17.265 -14.570 ;
      LAYER via ;
        RECT 17.075 6.880 17.335 7.140 ;
        RECT 17.075 6.560 17.335 6.820 ;
        RECT 17.075 6.240 17.335 6.500 ;
        RECT 17.075 5.920 17.335 6.180 ;
        RECT 17.075 5.600 17.335 5.860 ;
        RECT 17.075 5.280 17.335 5.540 ;
        RECT 17.075 4.960 17.335 5.220 ;
        RECT 17.075 4.640 17.335 4.900 ;
        RECT 17.075 4.320 17.335 4.580 ;
        RECT 17.075 4.000 17.335 4.260 ;
        RECT 17.075 3.680 17.335 3.940 ;
        RECT 17.075 3.360 17.335 3.620 ;
        RECT 17.075 3.040 17.335 3.300 ;
        RECT 17.075 2.720 17.335 2.980 ;
        RECT 17.075 2.400 17.335 2.660 ;
        RECT 17.075 2.080 17.335 2.340 ;
        RECT 14.855 -0.100 15.115 0.160 ;
        RECT 16.975 -9.720 17.235 -9.460 ;
        RECT 16.975 -10.040 17.235 -9.780 ;
        RECT 16.975 -10.360 17.235 -10.100 ;
        RECT 16.975 -10.680 17.235 -10.420 ;
        RECT 16.975 -11.000 17.235 -10.740 ;
        RECT 16.975 -11.320 17.235 -11.060 ;
        RECT 16.975 -11.640 17.235 -11.380 ;
        RECT 16.975 -11.960 17.235 -11.700 ;
        RECT 16.975 -12.280 17.235 -12.020 ;
        RECT 16.975 -12.600 17.235 -12.340 ;
        RECT 16.975 -12.920 17.235 -12.660 ;
        RECT 16.975 -13.240 17.235 -12.980 ;
        RECT 16.975 -13.560 17.235 -13.300 ;
        RECT 16.975 -13.880 17.235 -13.620 ;
        RECT 16.975 -14.200 17.235 -13.940 ;
        RECT 16.975 -14.520 17.235 -14.260 ;
        RECT 14.755 -16.700 15.015 -16.440 ;
      LAYER met2 ;
        RECT 17.045 1.995 17.365 7.345 ;
        RECT 14.775 -0.160 15.280 0.230 ;
        RECT 14.775 -16.370 15.180 -0.160 ;
        RECT 16.945 -14.605 17.265 -9.255 ;
        RECT 14.675 -16.760 15.280 -16.370 ;
    END
  END re_bl1
  PIN bl1
    ANTENNADIFFAREA 0.244800 ;
    PORT
      LAYER li1 ;
        RECT 18.705 5.340 20.045 5.590 ;
        RECT 18.605 -11.260 19.945 -11.010 ;
      LAYER mcon ;
        RECT 19.015 5.380 19.185 5.550 ;
        RECT 18.915 -11.220 19.085 -11.050 ;
      LAYER met1 ;
        RECT 18.395 7.655 19.235 8.215 ;
        RECT 18.975 5.590 19.235 7.655 ;
        RECT 18.955 5.320 19.245 5.590 ;
        RECT 15.425 0.610 15.700 0.830 ;
        RECT 18.975 0.610 19.235 5.320 ;
        RECT 15.425 0.405 19.235 0.610 ;
        RECT 18.295 -8.945 19.135 -8.385 ;
        RECT 18.875 -11.010 19.135 -8.945 ;
        RECT 18.855 -11.280 19.145 -11.010 ;
        RECT 15.325 -15.990 15.600 -15.770 ;
        RECT 18.875 -15.990 19.135 -11.280 ;
        RECT 15.325 -16.195 19.135 -15.990 ;
      LAYER via ;
        RECT 18.555 7.810 18.815 8.070 ;
        RECT 15.430 0.460 15.690 0.720 ;
        RECT 18.455 -8.790 18.715 -8.530 ;
        RECT 15.330 -16.140 15.590 -15.880 ;
      LAYER met2 ;
        RECT 18.395 8.210 18.965 8.220 ;
        RECT 17.570 7.930 18.965 8.210 ;
        RECT 18.395 7.645 18.965 7.930 ;
        RECT 15.420 -15.765 15.710 0.835 ;
        RECT 18.295 -8.390 18.865 -8.380 ;
        RECT 17.470 -8.670 18.865 -8.390 ;
        RECT 18.295 -8.955 18.865 -8.670 ;
        RECT 15.320 -16.190 15.710 -15.765 ;
    END
  END bl1
  PIN vdd
    ANTENNADIFFAREA 0.262800 ;
    PORT
      LAYER nwell ;
        RECT 18.255 2.305 19.235 5.590 ;
        RECT 18.155 -14.295 19.135 -11.010 ;
      LAYER li1 ;
        RECT 18.455 2.305 18.715 2.885 ;
        RECT 18.355 -14.295 18.615 -13.715 ;
      LAYER mcon ;
        RECT 18.505 2.450 18.675 2.620 ;
        RECT 18.405 -14.150 18.575 -13.980 ;
      LAYER met1 ;
        RECT 15.980 0.955 16.340 1.125 ;
        RECT 18.455 0.955 18.715 2.775 ;
        RECT 15.980 0.750 18.715 0.955 ;
        RECT 15.880 -15.645 16.240 -15.475 ;
        RECT 18.355 -15.645 18.615 -13.825 ;
        RECT 15.880 -15.850 18.615 -15.645 ;
      LAYER via ;
        RECT 16.025 0.815 16.285 1.075 ;
        RECT 15.925 -15.785 16.185 -15.525 ;
      LAYER met2 ;
        RECT 15.980 -15.470 16.345 1.130 ;
        RECT 15.880 -15.850 16.345 -15.470 ;
    END
    PORT
      LAYER nwell ;
        RECT -1.995 2.305 -1.015 5.590 ;
        RECT -2.095 -14.295 -1.115 -11.010 ;
      LAYER li1 ;
        RECT -1.795 2.305 -1.535 2.885 ;
        RECT -1.895 -14.295 -1.635 -13.715 ;
      LAYER mcon ;
        RECT -1.745 2.450 -1.575 2.620 ;
        RECT -1.845 -14.150 -1.675 -13.980 ;
      LAYER met1 ;
        RECT -4.270 0.955 -3.910 1.125 ;
        RECT -1.795 0.955 -1.535 2.775 ;
        RECT -4.270 0.750 -1.535 0.955 ;
        RECT -4.370 -15.645 -4.010 -15.475 ;
        RECT -1.895 -15.645 -1.635 -13.825 ;
        RECT -4.370 -15.850 -1.635 -15.645 ;
      LAYER via ;
        RECT -4.225 0.815 -3.965 1.075 ;
        RECT -4.325 -15.785 -4.065 -15.525 ;
      LAYER met2 ;
        RECT -4.270 -15.470 -3.905 1.130 ;
        RECT -4.370 -15.850 -3.905 -15.470 ;
    END
  END vdd
  PIN re_bl0
    ANTENNADIFFAREA 4.200000 ;
    PORT
      LAYER li1 ;
        RECT -3.160 1.990 -2.990 7.340 ;
        RECT -3.260 -14.610 -3.090 -9.260 ;
      LAYER mcon ;
        RECT -3.160 6.955 -2.990 7.125 ;
        RECT -3.160 6.595 -2.990 6.765 ;
        RECT -3.160 6.235 -2.990 6.405 ;
        RECT -3.160 5.875 -2.990 6.045 ;
        RECT -3.160 5.515 -2.990 5.685 ;
        RECT -3.160 5.155 -2.990 5.325 ;
        RECT -3.160 4.795 -2.990 4.965 ;
        RECT -3.160 4.435 -2.990 4.605 ;
        RECT -3.160 4.075 -2.990 4.245 ;
        RECT -3.160 3.715 -2.990 3.885 ;
        RECT -3.160 3.355 -2.990 3.525 ;
        RECT -3.160 2.995 -2.990 3.165 ;
        RECT -3.160 2.635 -2.990 2.805 ;
        RECT -3.160 2.275 -2.990 2.445 ;
        RECT -3.260 -9.645 -3.090 -9.475 ;
        RECT -3.260 -10.005 -3.090 -9.835 ;
        RECT -3.260 -10.365 -3.090 -10.195 ;
        RECT -3.260 -10.725 -3.090 -10.555 ;
        RECT -3.260 -11.085 -3.090 -10.915 ;
        RECT -3.260 -11.445 -3.090 -11.275 ;
        RECT -3.260 -11.805 -3.090 -11.635 ;
        RECT -3.260 -12.165 -3.090 -11.995 ;
        RECT -3.260 -12.525 -3.090 -12.355 ;
        RECT -3.260 -12.885 -3.090 -12.715 ;
        RECT -3.260 -13.245 -3.090 -13.075 ;
        RECT -3.260 -13.605 -3.090 -13.435 ;
        RECT -3.260 -13.965 -3.090 -13.795 ;
        RECT -3.260 -14.325 -3.090 -14.155 ;
      LAYER met1 ;
        RECT -3.205 2.345 -2.885 7.345 ;
        RECT -5.465 2.030 -2.885 2.345 ;
        RECT -5.465 -0.115 -5.100 2.030 ;
        RECT -3.205 1.990 -2.885 2.030 ;
        RECT -3.305 -14.255 -2.985 -9.255 ;
        RECT -5.565 -14.570 -2.985 -14.255 ;
        RECT -5.565 -16.715 -5.200 -14.570 ;
        RECT -3.305 -14.610 -2.985 -14.570 ;
      LAYER via ;
        RECT -3.175 6.880 -2.915 7.140 ;
        RECT -3.175 6.560 -2.915 6.820 ;
        RECT -3.175 6.240 -2.915 6.500 ;
        RECT -3.175 5.920 -2.915 6.180 ;
        RECT -3.175 5.600 -2.915 5.860 ;
        RECT -3.175 5.280 -2.915 5.540 ;
        RECT -3.175 4.960 -2.915 5.220 ;
        RECT -3.175 4.640 -2.915 4.900 ;
        RECT -3.175 4.320 -2.915 4.580 ;
        RECT -3.175 4.000 -2.915 4.260 ;
        RECT -3.175 3.680 -2.915 3.940 ;
        RECT -3.175 3.360 -2.915 3.620 ;
        RECT -3.175 3.040 -2.915 3.300 ;
        RECT -3.175 2.720 -2.915 2.980 ;
        RECT -3.175 2.400 -2.915 2.660 ;
        RECT -3.175 2.080 -2.915 2.340 ;
        RECT -5.395 -0.100 -5.135 0.160 ;
        RECT -3.275 -9.720 -3.015 -9.460 ;
        RECT -3.275 -10.040 -3.015 -9.780 ;
        RECT -3.275 -10.360 -3.015 -10.100 ;
        RECT -3.275 -10.680 -3.015 -10.420 ;
        RECT -3.275 -11.000 -3.015 -10.740 ;
        RECT -3.275 -11.320 -3.015 -11.060 ;
        RECT -3.275 -11.640 -3.015 -11.380 ;
        RECT -3.275 -11.960 -3.015 -11.700 ;
        RECT -3.275 -12.280 -3.015 -12.020 ;
        RECT -3.275 -12.600 -3.015 -12.340 ;
        RECT -3.275 -12.920 -3.015 -12.660 ;
        RECT -3.275 -13.240 -3.015 -12.980 ;
        RECT -3.275 -13.560 -3.015 -13.300 ;
        RECT -3.275 -13.880 -3.015 -13.620 ;
        RECT -3.275 -14.200 -3.015 -13.940 ;
        RECT -3.275 -14.520 -3.015 -14.260 ;
        RECT -5.495 -16.700 -5.235 -16.440 ;
      LAYER met2 ;
        RECT -3.205 1.995 -2.885 7.345 ;
        RECT -5.475 -0.160 -4.970 0.230 ;
        RECT -5.475 -16.370 -5.070 -0.160 ;
        RECT -3.305 -14.605 -2.985 -9.255 ;
        RECT -5.575 -16.760 -4.970 -16.370 ;
    END
  END re_bl0
  PIN bl0
    ANTENNADIFFAREA 0.244800 ;
    PORT
      LAYER li1 ;
        RECT -1.545 5.340 -0.205 5.590 ;
        RECT -1.645 -11.260 -0.305 -11.010 ;
      LAYER mcon ;
        RECT -1.235 5.380 -1.065 5.550 ;
        RECT -1.335 -11.220 -1.165 -11.050 ;
      LAYER met1 ;
        RECT -1.855 7.655 -1.015 8.215 ;
        RECT -1.275 5.590 -1.015 7.655 ;
        RECT -1.295 5.320 -1.005 5.590 ;
        RECT -4.825 0.610 -4.550 0.830 ;
        RECT -1.275 0.610 -1.015 5.320 ;
        RECT -4.825 0.405 -1.015 0.610 ;
        RECT -1.955 -8.945 -1.115 -8.385 ;
        RECT -1.375 -11.010 -1.115 -8.945 ;
        RECT -1.395 -11.280 -1.105 -11.010 ;
        RECT -4.925 -15.990 -4.650 -15.770 ;
        RECT -1.375 -15.990 -1.115 -11.280 ;
        RECT -4.925 -16.195 -1.115 -15.990 ;
      LAYER via ;
        RECT -1.695 7.810 -1.435 8.070 ;
        RECT -4.820 0.460 -4.560 0.720 ;
        RECT -1.795 -8.790 -1.535 -8.530 ;
        RECT -4.920 -16.140 -4.660 -15.880 ;
      LAYER met2 ;
        RECT -1.855 8.210 -1.285 8.220 ;
        RECT -2.680 7.930 -1.285 8.210 ;
        RECT -1.855 7.645 -1.285 7.930 ;
        RECT -4.830 -15.765 -4.540 0.835 ;
        RECT -1.955 -8.390 -1.385 -8.380 ;
        RECT -2.780 -8.670 -1.385 -8.390 ;
        RECT -1.955 -8.955 -1.385 -8.670 ;
        RECT -4.930 -16.190 -4.540 -15.765 ;
    END
  END bl0
  PIN br0
    ANTENNADIFFAREA 0.244800 ;
    PORT
      LAYER li1 ;
        RECT -1.545 3.190 -0.205 3.440 ;
        RECT -1.645 -13.410 -0.305 -13.160 ;
      LAYER mcon ;
        RECT -0.695 3.230 -0.525 3.400 ;
        RECT -0.795 -13.370 -0.625 -13.200 ;
      LAYER met1 ;
        RECT -0.755 7.650 0.135 8.230 ;
        RECT -0.755 5.590 -0.465 7.650 ;
        RECT -0.745 3.460 -0.485 5.590 ;
        RECT -0.755 3.190 -0.465 3.460 ;
        RECT -0.745 0.610 -0.485 3.190 ;
        RECT 2.950 0.610 3.225 0.830 ;
        RECT -0.745 0.405 3.225 0.610 ;
        RECT -0.745 0.400 -0.485 0.405 ;
        RECT -0.855 -8.950 0.035 -8.370 ;
        RECT -0.855 -11.010 -0.565 -8.950 ;
        RECT -0.845 -13.140 -0.585 -11.010 ;
        RECT -0.855 -13.410 -0.565 -13.140 ;
        RECT -0.845 -15.990 -0.585 -13.410 ;
        RECT 2.850 -15.990 3.125 -15.770 ;
        RECT -0.845 -16.195 3.125 -15.990 ;
        RECT -0.845 -16.200 -0.585 -16.195 ;
      LAYER via ;
        RECT -0.285 7.800 -0.025 8.060 ;
        RECT 2.955 0.460 3.215 0.720 ;
        RECT -0.385 -8.800 -0.125 -8.540 ;
        RECT 2.855 -16.140 3.115 -15.880 ;
      LAYER met2 ;
        RECT -0.460 7.960 1.275 8.230 ;
        RECT -0.460 7.655 0.130 7.960 ;
        RECT -0.560 -8.640 1.175 -8.370 ;
        RECT -0.560 -8.945 0.030 -8.640 ;
        RECT 2.945 -15.765 3.235 0.835 ;
        RECT 2.845 -16.190 3.235 -15.765 ;
    END
  END br0
  PIN re_br0
    ANTENNADIFFAREA 4.200000 ;
    PORT
      LAYER li1 ;
        RECT 1.115 1.990 1.285 7.340 ;
        RECT 1.015 -14.610 1.185 -9.260 ;
      LAYER mcon ;
        RECT 1.115 6.955 1.285 7.125 ;
        RECT 1.115 6.595 1.285 6.765 ;
        RECT 1.115 6.235 1.285 6.405 ;
        RECT 1.115 5.875 1.285 6.045 ;
        RECT 1.115 5.515 1.285 5.685 ;
        RECT 1.115 5.155 1.285 5.325 ;
        RECT 1.115 4.795 1.285 4.965 ;
        RECT 1.115 4.435 1.285 4.605 ;
        RECT 1.115 4.075 1.285 4.245 ;
        RECT 1.115 3.715 1.285 3.885 ;
        RECT 1.115 3.355 1.285 3.525 ;
        RECT 1.115 2.995 1.285 3.165 ;
        RECT 1.115 2.635 1.285 2.805 ;
        RECT 1.115 2.275 1.285 2.445 ;
        RECT 1.015 -9.645 1.185 -9.475 ;
        RECT 1.015 -10.005 1.185 -9.835 ;
        RECT 1.015 -10.365 1.185 -10.195 ;
        RECT 1.015 -10.725 1.185 -10.555 ;
        RECT 1.015 -11.085 1.185 -10.915 ;
        RECT 1.015 -11.445 1.185 -11.275 ;
        RECT 1.015 -11.805 1.185 -11.635 ;
        RECT 1.015 -12.165 1.185 -11.995 ;
        RECT 1.015 -12.525 1.185 -12.355 ;
        RECT 1.015 -12.885 1.185 -12.715 ;
        RECT 1.015 -13.245 1.185 -13.075 ;
        RECT 1.015 -13.605 1.185 -13.435 ;
        RECT 1.015 -13.965 1.185 -13.795 ;
        RECT 1.015 -14.325 1.185 -14.155 ;
      LAYER met1 ;
        RECT 1.070 1.730 1.390 7.345 ;
        RECT 1.070 1.525 3.985 1.730 ;
        RECT 3.705 -0.160 3.985 1.525 ;
        RECT 0.970 -14.870 1.290 -9.255 ;
        RECT 0.970 -15.075 3.885 -14.870 ;
        RECT 3.605 -16.760 3.885 -15.075 ;
      LAYER via ;
        RECT 1.100 6.880 1.360 7.140 ;
        RECT 1.100 6.560 1.360 6.820 ;
        RECT 1.100 6.240 1.360 6.500 ;
        RECT 1.100 5.920 1.360 6.180 ;
        RECT 1.100 5.600 1.360 5.860 ;
        RECT 1.100 5.280 1.360 5.540 ;
        RECT 1.100 4.960 1.360 5.220 ;
        RECT 1.100 4.640 1.360 4.900 ;
        RECT 1.100 4.320 1.360 4.580 ;
        RECT 1.100 4.000 1.360 4.260 ;
        RECT 1.100 3.680 1.360 3.940 ;
        RECT 1.100 3.360 1.360 3.620 ;
        RECT 1.100 3.040 1.360 3.300 ;
        RECT 1.100 2.720 1.360 2.980 ;
        RECT 1.100 2.400 1.360 2.660 ;
        RECT 1.100 2.080 1.360 2.340 ;
        RECT 3.710 -0.100 3.970 0.160 ;
        RECT 1.000 -9.720 1.260 -9.460 ;
        RECT 1.000 -10.040 1.260 -9.780 ;
        RECT 1.000 -10.360 1.260 -10.100 ;
        RECT 1.000 -10.680 1.260 -10.420 ;
        RECT 1.000 -11.000 1.260 -10.740 ;
        RECT 1.000 -11.320 1.260 -11.060 ;
        RECT 1.000 -11.640 1.260 -11.380 ;
        RECT 1.000 -11.960 1.260 -11.700 ;
        RECT 1.000 -12.280 1.260 -12.020 ;
        RECT 1.000 -12.600 1.260 -12.340 ;
        RECT 1.000 -12.920 1.260 -12.660 ;
        RECT 1.000 -13.240 1.260 -12.980 ;
        RECT 1.000 -13.560 1.260 -13.300 ;
        RECT 1.000 -13.880 1.260 -13.620 ;
        RECT 1.000 -14.200 1.260 -13.940 ;
        RECT 1.000 -14.520 1.260 -14.260 ;
        RECT 3.610 -16.700 3.870 -16.440 ;
      LAYER met2 ;
        RECT 1.070 1.995 1.390 7.345 ;
        RECT 0.970 -14.605 1.290 -9.255 ;
        RECT 3.480 -16.370 3.985 0.230 ;
        RECT 3.380 -16.760 3.985 -16.370 ;
    END
  END re_br0
  PIN VDD_HEADER0
    ANTENNAGATEAREA 0.108000 ;
    PORT
      LAYER li1 ;
        RECT -1.845 10.310 -1.285 10.595 ;
        RECT 18.405 10.310 18.965 10.595 ;
      LAYER mcon ;
        RECT -1.510 10.375 -1.340 10.545 ;
        RECT 18.740 10.375 18.910 10.545 ;
      LAYER met1 ;
        RECT -1.885 10.275 19.045 10.745 ;
      LAYER via ;
        RECT 5.665 10.365 5.925 10.625 ;
      LAYER met2 ;
        RECT 5.515 10.175 6.080 12.880 ;
    END
  END VDD_HEADER0
  PIN GND_HEADER0
    ANTENNAGATEAREA 0.054000 ;
    PORT
      LAYER li1 ;
        RECT -0.250 9.685 0.310 9.970 ;
      LAYER mcon ;
        RECT 0.085 9.750 0.255 9.920 ;
      LAYER met1 ;
        RECT -0.330 9.635 13.850 10.035 ;
      LAYER via ;
        RECT 7.790 9.695 8.050 9.955 ;
      LAYER met2 ;
        RECT 7.635 8.900 8.200 12.880 ;
    END
  END GND_HEADER0
  PIN VDD_HEADER1
    ANTENNAGATEAREA 0.108000 ;
    PORT
      LAYER li1 ;
        RECT -1.945 -6.290 -1.385 -6.005 ;
        RECT 18.305 -6.290 18.865 -6.005 ;
      LAYER mcon ;
        RECT -1.610 -6.225 -1.440 -6.055 ;
        RECT 18.640 -6.225 18.810 -6.055 ;
      LAYER met1 ;
        RECT -1.985 -6.005 18.715 -5.875 ;
        RECT -1.985 -6.290 18.940 -6.005 ;
        RECT -1.985 -6.345 18.715 -6.290 ;
      LAYER via ;
        RECT 10.065 -6.255 10.325 -5.995 ;
      LAYER met2 ;
        RECT 9.915 -6.445 10.480 12.880 ;
    END
  END VDD_HEADER1
  PIN GND_HEADER1
    ANTENNAGATEAREA 0.054000 ;
    PORT
      LAYER li1 ;
        RECT -0.350 -6.915 0.210 -6.630 ;
      LAYER mcon ;
        RECT -0.015 -6.850 0.155 -6.680 ;
      LAYER met1 ;
        RECT -0.430 -6.965 12.400 -6.565 ;
      LAYER via ;
        RECT 11.980 -6.890 12.240 -6.630 ;
      LAYER met2 ;
        RECT 11.835 -7.700 12.400 12.880 ;
    END
  END GND_HEADER1
  OBS
      LAYER nwell ;
        RECT -2.180 9.610 -1.180 10.640 ;
        RECT 18.070 9.610 19.070 10.640 ;
        RECT -1.935 9.555 -1.425 9.610 ;
      LAYER pwell ;
        RECT -0.590 8.980 0.420 9.600 ;
      LAYER nwell ;
        RECT 18.315 9.555 18.825 9.610 ;
      LAYER pwell ;
        RECT 19.660 8.980 20.670 9.600 ;
        RECT -3.330 0.215 -2.320 7.475 ;
        RECT -0.695 5.150 -0.075 5.720 ;
        RECT -0.725 4.650 -0.045 5.150 ;
        RECT -0.725 4.140 0.185 4.650 ;
        RECT -0.725 3.630 -0.045 4.140 ;
        RECT -0.695 3.060 -0.075 3.630 ;
        RECT 0.945 0.215 1.955 7.475 ;
        RECT 16.920 0.215 17.930 7.475 ;
        RECT 19.555 5.150 20.175 5.720 ;
        RECT 19.525 4.650 20.205 5.150 ;
        RECT 19.525 4.140 20.435 4.650 ;
        RECT 19.525 3.630 20.205 4.140 ;
        RECT 19.555 3.060 20.175 3.630 ;
        RECT 21.195 0.215 22.205 7.475 ;
      LAYER nwell ;
        RECT -2.280 -6.990 -1.280 -5.960 ;
        RECT 17.970 -6.990 18.970 -5.960 ;
        RECT -2.035 -7.045 -1.525 -6.990 ;
      LAYER pwell ;
        RECT -0.690 -7.620 0.320 -7.000 ;
      LAYER nwell ;
        RECT 18.215 -7.045 18.725 -6.990 ;
      LAYER pwell ;
        RECT 19.560 -7.620 20.570 -7.000 ;
        RECT -3.430 -16.385 -2.420 -9.125 ;
        RECT -0.795 -11.450 -0.175 -10.880 ;
        RECT -0.825 -11.950 -0.145 -11.450 ;
        RECT -0.825 -12.460 0.085 -11.950 ;
        RECT -0.825 -12.970 -0.145 -12.460 ;
        RECT -0.795 -13.540 -0.175 -12.970 ;
        RECT 0.845 -16.385 1.855 -9.125 ;
        RECT 16.820 -16.385 17.830 -9.125 ;
        RECT 19.455 -11.450 20.075 -10.880 ;
        RECT 19.425 -11.950 20.105 -11.450 ;
        RECT 19.425 -12.460 20.335 -11.950 ;
        RECT 19.425 -12.970 20.105 -12.460 ;
        RECT 19.455 -13.540 20.075 -12.970 ;
        RECT 21.095 -16.385 22.105 -9.125 ;
      LAYER li1 ;
        RECT -2.015 9.750 -1.845 10.080 ;
        RECT -1.515 9.750 -1.345 10.080 ;
        RECT 18.235 9.750 18.405 10.080 ;
        RECT 18.735 9.750 18.905 10.080 ;
        RECT 20.000 9.685 20.560 9.970 ;
        RECT -2.660 1.990 -2.490 7.340 ;
        RECT -1.860 5.925 -1.490 9.465 ;
        RECT -0.420 9.125 -0.250 9.455 ;
        RECT 0.080 9.125 0.250 9.455 ;
        RECT -0.240 5.925 0.110 8.790 ;
        RECT -1.535 5.060 -0.285 5.170 ;
        RECT -1.615 5.000 -0.205 5.060 ;
        RECT -1.615 4.730 -1.215 5.000 ;
        RECT -1.815 4.220 -1.565 4.550 ;
        RECT -1.385 4.400 -1.215 4.730 ;
        RECT -1.035 4.750 -0.705 4.830 ;
        RECT -1.035 4.580 -0.625 4.750 ;
        RECT -0.455 4.730 -0.205 5.000 ;
        RECT -0.795 4.560 -0.625 4.580 ;
        RECT -1.385 4.230 -1.025 4.400 ;
        RECT -0.795 4.390 -0.365 4.560 ;
        RECT -1.195 4.200 -1.025 4.230 ;
        RECT -1.615 3.780 -1.365 4.050 ;
        RECT -1.195 4.030 -0.705 4.200 ;
        RECT -1.035 3.950 -0.705 4.030 ;
        RECT -0.535 4.050 -0.365 4.390 ;
        RECT -0.195 4.230 0.055 4.560 ;
        RECT -0.535 3.780 -0.205 4.050 ;
        RECT -1.615 3.720 -0.205 3.780 ;
        RECT -1.535 3.610 -0.285 3.720 ;
        RECT 1.615 1.990 1.785 7.340 ;
        RECT 17.590 1.990 17.760 7.340 ;
        RECT 18.390 5.925 18.760 9.465 ;
        RECT 19.830 9.125 20.000 9.455 ;
        RECT 20.330 9.125 20.500 9.455 ;
        RECT 20.010 5.925 20.360 8.790 ;
        RECT 18.715 5.060 19.965 5.170 ;
        RECT 18.635 5.000 20.045 5.060 ;
        RECT 18.635 4.730 19.035 5.000 ;
        RECT 18.435 4.220 18.685 4.550 ;
        RECT 18.865 4.400 19.035 4.730 ;
        RECT 19.215 4.750 19.545 4.830 ;
        RECT 19.215 4.580 19.625 4.750 ;
        RECT 19.795 4.730 20.045 5.000 ;
        RECT 19.455 4.560 19.625 4.580 ;
        RECT 18.865 4.230 19.225 4.400 ;
        RECT 19.455 4.390 19.885 4.560 ;
        RECT 19.055 4.200 19.225 4.230 ;
        RECT 18.635 3.780 18.885 4.050 ;
        RECT 19.055 4.030 19.545 4.200 ;
        RECT 19.215 3.950 19.545 4.030 ;
        RECT 19.715 4.050 19.885 4.390 ;
        RECT 20.055 4.230 20.305 4.560 ;
        RECT 19.715 3.780 20.045 4.050 ;
        RECT 18.635 3.720 20.045 3.780 ;
        RECT 18.715 3.610 19.965 3.720 ;
        RECT 21.865 1.990 22.035 7.340 ;
        RECT -2.115 -6.850 -1.945 -6.520 ;
        RECT -1.615 -6.850 -1.445 -6.520 ;
        RECT 18.135 -6.850 18.305 -6.520 ;
        RECT 18.635 -6.850 18.805 -6.520 ;
        RECT 19.900 -6.915 20.460 -6.630 ;
        RECT -2.760 -14.610 -2.590 -9.260 ;
        RECT -1.960 -10.675 -1.590 -7.135 ;
        RECT -0.520 -7.475 -0.350 -7.145 ;
        RECT -0.020 -7.475 0.150 -7.145 ;
        RECT -0.340 -10.675 0.010 -7.810 ;
        RECT -1.635 -11.540 -0.385 -11.430 ;
        RECT -1.715 -11.600 -0.305 -11.540 ;
        RECT -1.715 -11.870 -1.315 -11.600 ;
        RECT -1.915 -12.380 -1.665 -12.050 ;
        RECT -1.485 -12.200 -1.315 -11.870 ;
        RECT -1.135 -11.850 -0.805 -11.770 ;
        RECT -1.135 -12.020 -0.725 -11.850 ;
        RECT -0.555 -11.870 -0.305 -11.600 ;
        RECT -0.895 -12.040 -0.725 -12.020 ;
        RECT -1.485 -12.370 -1.125 -12.200 ;
        RECT -0.895 -12.210 -0.465 -12.040 ;
        RECT -1.295 -12.400 -1.125 -12.370 ;
        RECT -1.715 -12.820 -1.465 -12.550 ;
        RECT -1.295 -12.570 -0.805 -12.400 ;
        RECT -1.135 -12.650 -0.805 -12.570 ;
        RECT -0.635 -12.550 -0.465 -12.210 ;
        RECT -0.295 -12.370 -0.045 -12.040 ;
        RECT -0.635 -12.820 -0.305 -12.550 ;
        RECT -1.715 -12.880 -0.305 -12.820 ;
        RECT -1.635 -12.990 -0.385 -12.880 ;
        RECT 1.515 -14.610 1.685 -9.260 ;
        RECT 17.490 -14.610 17.660 -9.260 ;
        RECT 18.290 -10.675 18.660 -7.135 ;
        RECT 19.730 -7.475 19.900 -7.145 ;
        RECT 20.230 -7.475 20.400 -7.145 ;
        RECT 19.910 -10.675 20.260 -7.810 ;
        RECT 18.615 -11.540 19.865 -11.430 ;
        RECT 18.535 -11.600 19.945 -11.540 ;
        RECT 18.535 -11.870 18.935 -11.600 ;
        RECT 18.335 -12.380 18.585 -12.050 ;
        RECT 18.765 -12.200 18.935 -11.870 ;
        RECT 19.115 -11.850 19.445 -11.770 ;
        RECT 19.115 -12.020 19.525 -11.850 ;
        RECT 19.695 -11.870 19.945 -11.600 ;
        RECT 19.355 -12.040 19.525 -12.020 ;
        RECT 18.765 -12.370 19.125 -12.200 ;
        RECT 19.355 -12.210 19.785 -12.040 ;
        RECT 18.955 -12.400 19.125 -12.370 ;
        RECT 18.535 -12.820 18.785 -12.550 ;
        RECT 18.955 -12.570 19.445 -12.400 ;
        RECT 19.115 -12.650 19.445 -12.570 ;
        RECT 19.615 -12.550 19.785 -12.210 ;
        RECT 19.955 -12.370 20.205 -12.040 ;
        RECT 19.615 -12.820 19.945 -12.550 ;
        RECT 18.535 -12.880 19.945 -12.820 ;
        RECT 18.615 -12.990 19.865 -12.880 ;
        RECT 21.765 -14.610 21.935 -9.260 ;
      LAYER mcon ;
        RECT -2.015 9.830 -1.845 10.000 ;
        RECT -1.515 9.830 -1.345 10.000 ;
        RECT 18.235 9.830 18.405 10.000 ;
        RECT 18.735 9.830 18.905 10.000 ;
        RECT 20.335 9.750 20.505 9.920 ;
        RECT -1.755 9.225 -1.585 9.395 ;
        RECT -2.660 6.950 -2.490 7.120 ;
        RECT -2.660 6.590 -2.490 6.760 ;
        RECT -2.660 6.230 -2.490 6.400 ;
        RECT -2.660 5.870 -2.490 6.040 ;
        RECT -0.420 9.205 -0.250 9.375 ;
        RECT 0.080 9.205 0.250 9.375 ;
        RECT 18.495 9.205 18.665 9.375 ;
        RECT -1.760 6.035 -1.590 6.205 ;
        RECT -0.160 8.570 0.010 8.740 ;
        RECT -0.175 6.030 -0.005 6.200 ;
        RECT 1.615 6.950 1.785 7.120 ;
        RECT 1.615 6.590 1.785 6.760 ;
        RECT 1.615 6.230 1.785 6.400 ;
        RECT -2.660 5.510 -2.490 5.680 ;
        RECT -2.660 5.150 -2.490 5.320 ;
        RECT 1.615 5.870 1.785 6.040 ;
        RECT 1.615 5.510 1.785 5.680 ;
        RECT 1.615 5.150 1.785 5.320 ;
        RECT -2.660 4.790 -2.490 4.960 ;
        RECT -2.660 4.430 -2.490 4.600 ;
        RECT -2.660 4.070 -2.490 4.240 ;
        RECT -1.735 4.300 -1.565 4.470 ;
        RECT 1.615 4.790 1.785 4.960 ;
        RECT -2.660 3.710 -2.490 3.880 ;
        RECT -0.195 4.310 -0.025 4.480 ;
        RECT 1.615 4.430 1.785 4.600 ;
        RECT 1.615 4.070 1.785 4.240 ;
        RECT 1.615 3.710 1.785 3.880 ;
        RECT -2.660 3.350 -2.490 3.520 ;
        RECT -2.660 2.990 -2.490 3.160 ;
        RECT -2.660 2.630 -2.490 2.800 ;
        RECT -2.660 2.270 -2.490 2.440 ;
        RECT 1.615 3.350 1.785 3.520 ;
        RECT 1.615 2.990 1.785 3.160 ;
        RECT 1.615 2.630 1.785 2.800 ;
        RECT 1.615 2.270 1.785 2.440 ;
        RECT 17.590 6.950 17.760 7.120 ;
        RECT 17.590 6.590 17.760 6.760 ;
        RECT 17.590 6.230 17.760 6.400 ;
        RECT 17.590 5.870 17.760 6.040 ;
        RECT 19.830 9.205 20.000 9.375 ;
        RECT 20.330 9.205 20.500 9.375 ;
        RECT 18.490 6.035 18.660 6.205 ;
        RECT 20.090 8.565 20.260 8.735 ;
        RECT 20.075 6.030 20.245 6.200 ;
        RECT 21.865 6.950 22.035 7.120 ;
        RECT 21.865 6.590 22.035 6.760 ;
        RECT 21.865 6.230 22.035 6.400 ;
        RECT 17.590 5.510 17.760 5.680 ;
        RECT 17.590 5.150 17.760 5.320 ;
        RECT 21.865 5.870 22.035 6.040 ;
        RECT 21.865 5.510 22.035 5.680 ;
        RECT 21.865 5.150 22.035 5.320 ;
        RECT 17.590 4.790 17.760 4.960 ;
        RECT 17.590 4.430 17.760 4.600 ;
        RECT 17.590 4.070 17.760 4.240 ;
        RECT 18.515 4.300 18.685 4.470 ;
        RECT 21.865 4.790 22.035 4.960 ;
        RECT 17.590 3.710 17.760 3.880 ;
        RECT 20.055 4.310 20.225 4.480 ;
        RECT 21.865 4.430 22.035 4.600 ;
        RECT 21.865 4.070 22.035 4.240 ;
        RECT 21.865 3.710 22.035 3.880 ;
        RECT 17.590 3.350 17.760 3.520 ;
        RECT 17.590 2.990 17.760 3.160 ;
        RECT 17.590 2.630 17.760 2.800 ;
        RECT 17.590 2.270 17.760 2.440 ;
        RECT 21.865 3.350 22.035 3.520 ;
        RECT 21.865 2.990 22.035 3.160 ;
        RECT 21.865 2.630 22.035 2.800 ;
        RECT 21.865 2.270 22.035 2.440 ;
        RECT -2.115 -6.770 -1.945 -6.600 ;
        RECT -1.615 -6.770 -1.445 -6.600 ;
        RECT 18.135 -6.770 18.305 -6.600 ;
        RECT 18.635 -6.770 18.805 -6.600 ;
        RECT 20.235 -6.850 20.405 -6.680 ;
        RECT -1.855 -7.375 -1.685 -7.205 ;
        RECT -2.760 -9.650 -2.590 -9.480 ;
        RECT -2.760 -10.010 -2.590 -9.840 ;
        RECT -2.760 -10.370 -2.590 -10.200 ;
        RECT -2.760 -10.730 -2.590 -10.560 ;
        RECT -0.520 -7.395 -0.350 -7.225 ;
        RECT -0.020 -7.395 0.150 -7.225 ;
        RECT 18.395 -7.380 18.565 -7.210 ;
        RECT -1.860 -10.565 -1.690 -10.395 ;
        RECT -0.260 -8.030 -0.090 -7.860 ;
        RECT -0.275 -10.570 -0.105 -10.400 ;
        RECT 1.515 -9.650 1.685 -9.480 ;
        RECT 1.515 -10.010 1.685 -9.840 ;
        RECT 1.515 -10.370 1.685 -10.200 ;
        RECT -2.760 -11.090 -2.590 -10.920 ;
        RECT -2.760 -11.450 -2.590 -11.280 ;
        RECT 1.515 -10.730 1.685 -10.560 ;
        RECT 1.515 -11.090 1.685 -10.920 ;
        RECT 1.515 -11.450 1.685 -11.280 ;
        RECT -2.760 -11.810 -2.590 -11.640 ;
        RECT -2.760 -12.170 -2.590 -12.000 ;
        RECT -2.760 -12.530 -2.590 -12.360 ;
        RECT -1.835 -12.300 -1.665 -12.130 ;
        RECT 1.515 -11.810 1.685 -11.640 ;
        RECT -2.760 -12.890 -2.590 -12.720 ;
        RECT -0.295 -12.290 -0.125 -12.120 ;
        RECT 1.515 -12.170 1.685 -12.000 ;
        RECT 1.515 -12.530 1.685 -12.360 ;
        RECT 1.515 -12.890 1.685 -12.720 ;
        RECT -2.760 -13.250 -2.590 -13.080 ;
        RECT -2.760 -13.610 -2.590 -13.440 ;
        RECT -2.760 -13.970 -2.590 -13.800 ;
        RECT -2.760 -14.330 -2.590 -14.160 ;
        RECT 1.515 -13.250 1.685 -13.080 ;
        RECT 1.515 -13.610 1.685 -13.440 ;
        RECT 1.515 -13.970 1.685 -13.800 ;
        RECT 1.515 -14.330 1.685 -14.160 ;
        RECT 17.490 -9.650 17.660 -9.480 ;
        RECT 17.490 -10.010 17.660 -9.840 ;
        RECT 17.490 -10.370 17.660 -10.200 ;
        RECT 17.490 -10.730 17.660 -10.560 ;
        RECT 19.730 -7.395 19.900 -7.225 ;
        RECT 20.230 -7.395 20.400 -7.225 ;
        RECT 18.390 -10.565 18.560 -10.395 ;
        RECT 19.990 -8.030 20.160 -7.860 ;
        RECT 19.975 -10.570 20.145 -10.400 ;
        RECT 21.765 -9.650 21.935 -9.480 ;
        RECT 21.765 -10.010 21.935 -9.840 ;
        RECT 21.765 -10.370 21.935 -10.200 ;
        RECT 17.490 -11.090 17.660 -10.920 ;
        RECT 17.490 -11.450 17.660 -11.280 ;
        RECT 21.765 -10.730 21.935 -10.560 ;
        RECT 21.765 -11.090 21.935 -10.920 ;
        RECT 21.765 -11.450 21.935 -11.280 ;
        RECT 17.490 -11.810 17.660 -11.640 ;
        RECT 17.490 -12.170 17.660 -12.000 ;
        RECT 17.490 -12.530 17.660 -12.360 ;
        RECT 18.415 -12.300 18.585 -12.130 ;
        RECT 21.765 -11.810 21.935 -11.640 ;
        RECT 17.490 -12.890 17.660 -12.720 ;
        RECT 19.955 -12.290 20.125 -12.120 ;
        RECT 21.765 -12.170 21.935 -12.000 ;
        RECT 21.765 -12.530 21.935 -12.360 ;
        RECT 21.765 -12.890 21.935 -12.720 ;
        RECT 17.490 -13.250 17.660 -13.080 ;
        RECT 17.490 -13.610 17.660 -13.440 ;
        RECT 17.490 -13.970 17.660 -13.800 ;
        RECT 17.490 -14.330 17.660 -14.160 ;
        RECT 21.765 -13.250 21.935 -13.080 ;
        RECT 21.765 -13.610 21.935 -13.440 ;
        RECT 21.765 -13.970 21.935 -13.800 ;
        RECT 21.765 -14.330 21.935 -14.160 ;
      LAYER met1 ;
        RECT -2.060 9.745 -1.740 10.065 ;
        RECT -1.545 9.770 -1.315 10.080 ;
        RECT -1.500 9.605 -1.360 9.770 ;
        RECT 18.190 9.745 18.510 10.065 ;
        RECT 18.705 9.770 18.935 10.080 ;
        RECT 18.750 9.605 18.890 9.770 ;
        RECT 20.200 9.685 20.635 9.970 ;
        RECT -1.755 9.465 -1.360 9.605 ;
        RECT 18.495 9.465 18.890 9.605 ;
        RECT -1.860 9.075 -1.490 9.465 ;
        RECT -0.495 9.120 -0.145 9.455 ;
        RECT 0.050 9.145 0.280 9.455 ;
        RECT 0.095 8.980 0.235 9.145 ;
        RECT 18.390 9.085 18.760 9.465 ;
        RECT 19.755 9.120 20.105 9.455 ;
        RECT 20.300 9.145 20.530 9.455 ;
        RECT 20.345 8.980 20.485 9.145 ;
        RECT -0.160 8.840 0.235 8.980 ;
        RECT 20.090 8.840 20.485 8.980 ;
        RECT -0.240 8.480 0.110 8.840 ;
        RECT 20.010 8.480 20.360 8.840 ;
        RECT -3.000 7.940 -2.680 8.200 ;
        RECT 1.275 7.940 1.595 8.200 ;
        RECT 17.250 7.940 17.570 8.200 ;
        RECT 21.525 7.940 21.845 8.200 ;
        RECT -2.900 7.625 -2.740 7.940 ;
        RECT 1.375 7.625 1.535 7.940 ;
        RECT 17.350 7.625 17.510 7.940 ;
        RECT 21.625 7.625 21.785 7.940 ;
        RECT -2.900 7.485 -2.505 7.625 ;
        RECT 1.375 7.485 1.770 7.625 ;
        RECT 17.350 7.485 17.745 7.625 ;
        RECT 21.625 7.485 22.020 7.625 ;
        RECT -2.645 7.320 -2.505 7.485 ;
        RECT 1.630 7.320 1.770 7.485 ;
        RECT 17.605 7.320 17.745 7.485 ;
        RECT 21.880 7.320 22.020 7.485 ;
        RECT -2.690 1.990 -2.460 7.320 ;
        RECT -1.795 5.170 -1.535 6.300 ;
        RECT -0.205 5.590 0.035 6.300 ;
        RECT -1.795 4.850 -1.475 5.170 ;
        RECT -1.795 4.530 -1.535 4.850 ;
        RECT -0.225 4.550 0.035 5.590 ;
        RECT -1.795 4.240 -1.505 4.530 ;
        RECT -1.795 3.190 -1.535 4.240 ;
        RECT -0.285 4.230 0.035 4.550 ;
        RECT -0.225 3.190 0.035 4.230 ;
        RECT 1.585 1.990 1.815 7.320 ;
        RECT 17.560 1.990 17.790 7.320 ;
        RECT 18.455 5.170 18.715 6.300 ;
        RECT 20.045 5.590 20.285 6.300 ;
        RECT 18.455 4.850 18.775 5.170 ;
        RECT 18.455 4.530 18.715 4.850 ;
        RECT 20.025 4.550 20.285 5.590 ;
        RECT 18.455 4.240 18.745 4.530 ;
        RECT 18.455 3.190 18.715 4.240 ;
        RECT 19.965 4.230 20.285 4.550 ;
        RECT 20.025 3.190 20.285 4.230 ;
        RECT 21.835 1.990 22.065 7.320 ;
        RECT -2.160 -6.855 -1.840 -6.535 ;
        RECT -1.645 -6.830 -1.415 -6.520 ;
        RECT -1.600 -6.995 -1.460 -6.830 ;
        RECT 18.090 -6.855 18.410 -6.535 ;
        RECT 18.605 -6.830 18.835 -6.520 ;
        RECT 18.650 -6.995 18.790 -6.830 ;
        RECT 20.100 -6.915 20.535 -6.630 ;
        RECT -1.855 -7.135 -1.460 -6.995 ;
        RECT 18.395 -7.135 18.790 -6.995 ;
        RECT -1.960 -7.485 -1.590 -7.135 ;
        RECT -0.595 -7.480 -0.245 -7.145 ;
        RECT -0.050 -7.455 0.180 -7.145 ;
        RECT -0.005 -7.620 0.135 -7.455 ;
        RECT 18.290 -7.465 18.660 -7.135 ;
        RECT 19.655 -7.480 20.005 -7.145 ;
        RECT 20.200 -7.455 20.430 -7.145 ;
        RECT 20.245 -7.620 20.385 -7.455 ;
        RECT -0.260 -7.760 0.135 -7.620 ;
        RECT 19.990 -7.760 20.385 -7.620 ;
        RECT -0.340 -8.175 0.010 -7.760 ;
        RECT 19.910 -8.110 20.260 -7.760 ;
        RECT -3.100 -8.660 -2.780 -8.400 ;
        RECT 1.175 -8.660 1.495 -8.400 ;
        RECT 17.150 -8.660 17.470 -8.400 ;
        RECT 21.425 -8.660 21.745 -8.400 ;
        RECT -3.000 -8.975 -2.840 -8.660 ;
        RECT 1.275 -8.975 1.435 -8.660 ;
        RECT 17.250 -8.975 17.410 -8.660 ;
        RECT 21.525 -8.975 21.685 -8.660 ;
        RECT -3.000 -9.115 -2.605 -8.975 ;
        RECT 1.275 -9.115 1.670 -8.975 ;
        RECT 17.250 -9.115 17.645 -8.975 ;
        RECT 21.525 -9.115 21.920 -8.975 ;
        RECT -2.745 -9.280 -2.605 -9.115 ;
        RECT 1.530 -9.280 1.670 -9.115 ;
        RECT 17.505 -9.280 17.645 -9.115 ;
        RECT 21.780 -9.280 21.920 -9.115 ;
        RECT -2.790 -14.610 -2.560 -9.280 ;
        RECT -1.895 -11.430 -1.635 -10.300 ;
        RECT -0.305 -11.010 -0.065 -10.300 ;
        RECT -1.895 -11.750 -1.575 -11.430 ;
        RECT -1.895 -12.070 -1.635 -11.750 ;
        RECT -0.325 -12.050 -0.065 -11.010 ;
        RECT -1.895 -12.360 -1.605 -12.070 ;
        RECT -1.895 -13.410 -1.635 -12.360 ;
        RECT -0.385 -12.370 -0.065 -12.050 ;
        RECT -0.325 -13.410 -0.065 -12.370 ;
        RECT 1.485 -14.610 1.715 -9.280 ;
        RECT 17.460 -14.610 17.690 -9.280 ;
        RECT 18.355 -11.430 18.615 -10.300 ;
        RECT 19.945 -11.010 20.185 -10.300 ;
        RECT 18.355 -11.750 18.675 -11.430 ;
        RECT 18.355 -12.070 18.615 -11.750 ;
        RECT 19.925 -12.050 20.185 -11.010 ;
        RECT 18.355 -12.360 18.645 -12.070 ;
        RECT 18.355 -13.410 18.615 -12.360 ;
        RECT 19.865 -12.370 20.185 -12.050 ;
        RECT 19.925 -13.410 20.185 -12.370 ;
        RECT 21.735 -14.610 21.965 -9.280 ;
      LAYER via ;
        RECT -1.765 4.880 -1.505 5.140 ;
        RECT -0.255 4.260 0.005 4.520 ;
        RECT 18.485 4.880 18.745 5.140 ;
        RECT 19.995 4.260 20.255 4.520 ;
        RECT -1.865 -11.720 -1.605 -11.460 ;
        RECT -0.355 -12.340 -0.095 -12.080 ;
        RECT 18.385 -11.720 18.645 -11.460 ;
        RECT 19.895 -12.340 20.155 -12.080 ;
      LAYER met2 ;
        RECT -1.815 4.850 0.055 5.170 ;
        RECT 18.435 4.850 20.305 5.170 ;
        RECT -1.815 4.230 0.055 4.550 ;
        RECT 18.435 4.230 20.305 4.550 ;
        RECT -1.815 3.610 0.055 3.930 ;
        RECT 18.435 3.610 20.305 3.930 ;
        RECT -1.915 -11.750 -0.045 -11.430 ;
        RECT 18.335 -11.750 20.205 -11.430 ;
        RECT -1.915 -12.370 -0.045 -12.050 ;
        RECT 18.335 -12.370 20.205 -12.050 ;
        RECT -1.915 -12.990 -0.045 -12.670 ;
        RECT 18.335 -12.990 20.205 -12.670 ;
  END
END array
MACRO 1T1R_300U
  CLASS BLOCK ;
  FOREIGN 1T1R_300U ;
  ORIGIN 0.920 9.900 ;
  SIZE 1.010 BY 4.365 ;
  PIN G
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER li1 ;
        RECT -0.585 -9.900 -0.025 -9.615 ;
      LAYER mcon ;
        RECT -0.250 -9.850 -0.080 -9.680 ;
      LAYER met1 ;
        RECT -0.385 -9.900 0.050 -9.615 ;
      LAYER via ;
        RECT -0.300 -9.875 -0.040 -9.615 ;
      LAYER met2 ;
        RECT -0.385 -9.875 0.050 -9.615 ;
    END
  END G
  PIN S
    ANTENNADIFFAREA 0.900000 ;
    PORT
      LAYER li1 ;
        RECT -0.750 -9.440 -0.580 -6.455 ;
      LAYER mcon ;
        RECT -0.750 -7.005 -0.580 -6.835 ;
        RECT -0.750 -7.365 -0.580 -7.195 ;
        RECT -0.750 -7.725 -0.580 -7.555 ;
        RECT -0.750 -8.085 -0.580 -7.915 ;
        RECT -0.750 -8.445 -0.580 -8.275 ;
        RECT -0.750 -8.805 -0.580 -8.635 ;
        RECT -0.750 -9.165 -0.580 -8.995 ;
      LAYER met1 ;
        RECT -0.795 -9.440 -0.475 -6.450 ;
      LAYER via ;
        RECT -0.765 -6.995 -0.505 -6.735 ;
        RECT -0.765 -7.315 -0.505 -7.055 ;
        RECT -0.765 -7.635 -0.505 -7.375 ;
        RECT -0.765 -7.955 -0.505 -7.695 ;
        RECT -0.765 -8.275 -0.505 -8.015 ;
        RECT -0.765 -8.595 -0.505 -8.335 ;
        RECT -0.765 -8.915 -0.505 -8.655 ;
        RECT -0.765 -9.235 -0.505 -8.975 ;
      LAYER met2 ;
        RECT -0.795 -9.370 -0.475 -6.450 ;
    END
  END S
  OBS
      LAYER pwell ;
        RECT -0.920 -9.570 0.090 -6.310 ;
      LAYER li1 ;
        RECT -0.250 -9.440 -0.080 -6.455 ;
      LAYER mcon ;
        RECT -0.250 -7.005 -0.080 -6.835 ;
        RECT -0.250 -7.365 -0.080 -7.195 ;
        RECT -0.250 -7.725 -0.080 -7.555 ;
        RECT -0.250 -8.085 -0.080 -7.915 ;
        RECT -0.250 -8.445 -0.080 -8.275 ;
        RECT -0.250 -8.805 -0.080 -8.635 ;
        RECT -0.250 -9.165 -0.080 -8.995 ;
      LAYER met1 ;
        RECT -0.590 -5.855 -0.270 -5.595 ;
        RECT -0.490 -6.170 -0.330 -5.855 ;
        RECT -0.490 -6.310 -0.095 -6.170 ;
        RECT -0.235 -6.475 -0.095 -6.310 ;
        RECT -0.280 -9.440 -0.050 -6.475 ;
  END
END 1T1R_300U
MACRO 1T1R_100U
  CLASS BLOCK ;
  FOREIGN 1T1R_100U ;
  ORIGIN 0.920 8.065 ;
  SIZE 1.010 BY 2.530 ;
  PIN G
    ANTENNAGATEAREA 0.150000 ;
    PORT
      LAYER li1 ;
        RECT -0.580 -8.065 -0.020 -7.780 ;
      LAYER mcon ;
        RECT -0.245 -8.015 -0.075 -7.845 ;
      LAYER met1 ;
        RECT -0.380 -8.065 0.055 -7.780 ;
      LAYER via ;
        RECT -0.295 -8.040 -0.035 -7.780 ;
      LAYER met2 ;
        RECT -0.380 -8.040 0.055 -7.780 ;
    END
  END G
  PIN S
    ANTENNADIFFAREA 0.300000 ;
    PORT
      LAYER li1 ;
        RECT -0.750 -7.405 -0.580 -6.455 ;
      LAYER mcon ;
        RECT -0.750 -6.825 -0.580 -6.655 ;
        RECT -0.750 -7.185 -0.580 -7.015 ;
      LAYER met1 ;
        RECT -0.795 -7.410 -0.475 -6.450 ;
      LAYER via ;
        RECT -0.765 -6.890 -0.505 -6.630 ;
        RECT -0.765 -7.210 -0.505 -6.950 ;
      LAYER met2 ;
        RECT -0.795 -7.640 -0.475 -6.450 ;
    END
  END S
  OBS
      LAYER pwell ;
        RECT -0.920 -7.570 0.090 -6.310 ;
      LAYER li1 ;
        RECT -0.250 -7.405 -0.080 -6.455 ;
      LAYER mcon ;
        RECT -0.250 -6.830 -0.080 -6.660 ;
        RECT -0.250 -7.190 -0.080 -7.020 ;
      LAYER met1 ;
        RECT -0.590 -5.855 -0.270 -5.595 ;
        RECT -0.490 -6.170 -0.330 -5.855 ;
        RECT -0.490 -6.310 -0.095 -6.170 ;
        RECT -0.235 -6.475 -0.095 -6.310 ;
        RECT -0.280 -7.410 -0.050 -6.475 ;
  END
END 1T1R_100U
MACRO 1T1R_036U
  CLASS BLOCK ;
  FOREIGN 1T1R_036U ;
  ORIGIN 0.915 6.930 ;
  SIZE 1.000 BY 0.620 ;
  PIN G
    ANTENNAGATEAREA 0.054000 ;
    PORT
      LAYER li1 ;
        RECT -0.580 -7.300 -0.020 -7.015 ;
      LAYER mcon ;
        RECT -0.245 -7.250 -0.075 -7.080 ;
      LAYER met1 ;
        RECT -0.380 -7.300 0.055 -7.015 ;
      LAYER via ;
        RECT -0.295 -7.275 -0.035 -7.015 ;
      LAYER met2 ;
        RECT -0.380 -7.275 0.055 -7.015 ;
    END
  END G
  PIN S
    ANTENNADIFFAREA 0.108000 ;
    PORT
      LAYER li1 ;
        RECT -0.750 -6.785 -0.580 -6.455 ;
      LAYER mcon ;
        RECT -0.750 -6.705 -0.580 -6.535 ;
      LAYER met1 ;
        RECT -0.795 -6.770 -0.475 -6.450 ;
      LAYER via ;
        RECT -0.765 -6.740 -0.505 -6.480 ;
      LAYER met2 ;
        RECT -0.795 -6.770 -0.475 -6.450 ;
    END
  END S
  OBS
      LAYER pwell ;
        RECT -0.920 -6.930 0.090 -6.310 ;
      LAYER li1 ;
        RECT -0.250 -6.785 -0.080 -6.455 ;
      LAYER mcon ;
        RECT -0.250 -6.705 -0.080 -6.535 ;
      LAYER met1 ;
        RECT -0.590 -5.855 -0.270 -5.595 ;
        RECT -0.490 -6.170 -0.330 -5.855 ;
        RECT -0.490 -6.310 -0.095 -6.170 ;
        RECT -0.235 -6.475 -0.095 -6.310 ;
        RECT -0.280 -6.785 -0.050 -6.475 ;
  END
END 1T1R_036U
MACRO RRAM
  CLASS BLOCK ;
  FOREIGN RRAM ;
  ORIGIN 4.075 -9.735 ;
  SIZE 0.380 BY 0.380 ;
  PIN BE
    PORT
      LAYER met1 ;
        RECT -4.045 9.795 -3.725 10.055 ;
    END
  END BE
END RRAM
MACRO rram_test
  CLASS BLOCK ;
  FOREIGN rram_test ;
  ORIGIN 18.240 72.000 ;
  SIZE 65.120 BY 237.250 ;
  PIN p1T1R_WL
    ANTENNAGATEAREA 1.704000 ;
    PORT
      LAYER li1 ;
        RECT -4.520 1.505 -3.960 1.790 ;
        RECT -3.305 0.740 -2.745 1.025 ;
        RECT -2.255 -1.095 -1.695 -0.810 ;
        RECT -1.205 -5.105 -0.850 -4.820 ;
      LAYER mcon ;
        RECT -4.185 1.555 -4.015 1.725 ;
        RECT -2.970 0.790 -2.800 0.960 ;
        RECT -1.920 -1.045 -1.750 -0.875 ;
        RECT -1.115 -5.025 -0.945 -4.855 ;
      LAYER met1 ;
        RECT -4.320 1.025 -3.885 1.790 ;
        RECT -4.320 0.740 -2.670 1.025 ;
        RECT -4.320 -0.810 -3.885 0.740 ;
        RECT -4.320 -1.055 -1.620 -0.810 ;
        RECT -2.055 -4.655 -1.620 -1.055 ;
        RECT -2.055 -5.225 -0.695 -4.655 ;
      LAYER via ;
        RECT -4.235 1.530 -3.975 1.790 ;
        RECT -3.020 0.765 -2.760 1.025 ;
        RECT -1.970 -1.070 -1.710 -0.810 ;
        RECT -1.165 -5.065 -0.905 -4.805 ;
      LAYER met2 ;
        RECT -12.375 5.570 -10.560 7.350 ;
        RECT -11.010 1.790 -10.705 5.570 ;
        RECT -11.010 1.530 -3.885 1.790 ;
        RECT -3.105 0.765 -2.670 1.025 ;
        RECT -2.055 -1.070 -1.620 -0.810 ;
        RECT -1.350 -5.230 -0.690 -4.655 ;
    END
  END p1T1R_WL
  PIN p036_SL
    ANTENNADIFFAREA 0.108000 ;
    PORT
      LAYER li1 ;
        RECT -4.690 2.020 -4.520 2.350 ;
      LAYER mcon ;
        RECT -4.690 2.100 -4.520 2.270 ;
      LAYER met1 ;
        RECT -4.735 2.035 -4.415 2.355 ;
      LAYER via ;
        RECT -4.705 2.065 -4.445 2.325 ;
      LAYER met2 ;
        RECT -10.420 5.570 -8.605 7.350 ;
        RECT -9.110 2.355 -8.810 5.570 ;
        RECT -9.110 2.035 -4.415 2.355 ;
    END
  END p036_SL
  PIN p700_SL
    ANTENNADIFFAREA 2.100000 ;
    PORT
      LAYER li1 ;
        RECT -1.385 -3.000 -1.215 2.350 ;
      LAYER mcon ;
        RECT -1.385 1.965 -1.215 2.135 ;
        RECT -1.385 1.605 -1.215 1.775 ;
        RECT -1.385 1.245 -1.215 1.415 ;
        RECT -1.385 0.885 -1.215 1.055 ;
        RECT -1.385 0.525 -1.215 0.695 ;
        RECT -1.385 0.165 -1.215 0.335 ;
        RECT -1.385 -0.195 -1.215 -0.025 ;
        RECT -1.385 -0.555 -1.215 -0.385 ;
        RECT -1.385 -0.915 -1.215 -0.745 ;
        RECT -1.385 -1.275 -1.215 -1.105 ;
        RECT -1.385 -1.635 -1.215 -1.465 ;
        RECT -1.385 -1.995 -1.215 -1.825 ;
        RECT -1.385 -2.355 -1.215 -2.185 ;
        RECT -1.385 -2.715 -1.215 -2.545 ;
      LAYER met1 ;
        RECT -1.430 -3.000 -1.110 2.355 ;
      LAYER via ;
        RECT -1.400 1.890 -1.140 2.150 ;
        RECT -1.400 1.570 -1.140 1.830 ;
        RECT -1.400 1.250 -1.140 1.510 ;
        RECT -1.400 0.930 -1.140 1.190 ;
        RECT -1.400 0.610 -1.140 0.870 ;
        RECT -1.400 0.290 -1.140 0.550 ;
        RECT -1.400 -0.030 -1.140 0.230 ;
        RECT -1.400 -0.350 -1.140 -0.090 ;
        RECT -1.400 -0.670 -1.140 -0.410 ;
        RECT -1.400 -0.990 -1.140 -0.730 ;
        RECT -1.400 -1.310 -1.140 -1.050 ;
        RECT -1.400 -1.630 -1.140 -1.370 ;
        RECT -1.400 -1.950 -1.140 -1.690 ;
        RECT -1.400 -2.270 -1.140 -2.010 ;
        RECT -1.400 -2.590 -1.140 -2.330 ;
        RECT -1.400 -2.910 -1.140 -2.650 ;
      LAYER met2 ;
        RECT -18.240 5.570 -16.425 7.350 ;
        RECT -17.045 -2.310 -16.570 5.570 ;
        RECT -1.430 -2.310 -1.110 2.355 ;
        RECT -17.045 -2.600 -1.110 -2.310 ;
        RECT -1.430 -2.995 -1.110 -2.600 ;
    END
  END p700_SL
  PIN p300_SL
    ANTENNADIFFAREA 0.900000 ;
    PORT
      LAYER li1 ;
        RECT -2.420 -0.635 -2.250 2.350 ;
      LAYER mcon ;
        RECT -2.420 1.800 -2.250 1.970 ;
        RECT -2.420 1.440 -2.250 1.610 ;
        RECT -2.420 1.080 -2.250 1.250 ;
        RECT -2.420 0.720 -2.250 0.890 ;
        RECT -2.420 0.360 -2.250 0.530 ;
        RECT -2.420 0.000 -2.250 0.170 ;
        RECT -2.420 -0.360 -2.250 -0.190 ;
      LAYER met1 ;
        RECT -2.465 -0.635 -2.145 2.355 ;
      LAYER via ;
        RECT -2.435 1.810 -2.175 2.070 ;
        RECT -2.435 1.490 -2.175 1.750 ;
        RECT -2.435 1.170 -2.175 1.430 ;
        RECT -2.435 0.850 -2.175 1.110 ;
        RECT -2.435 0.530 -2.175 0.790 ;
        RECT -2.435 0.210 -2.175 0.470 ;
        RECT -2.435 -0.110 -2.175 0.150 ;
        RECT -2.435 -0.430 -2.175 -0.170 ;
      LAYER met2 ;
        RECT -16.285 5.570 -14.470 7.350 ;
        RECT -15.090 -0.175 -14.615 5.570 ;
        RECT -2.465 -0.175 -2.145 2.355 ;
        RECT -15.090 -0.435 -2.145 -0.175 ;
        RECT -2.465 -0.565 -2.145 -0.435 ;
    END
  END p300_SL
  PIN p100_SL
    ANTENNADIFFAREA 0.300000 ;
    PORT
      LAYER li1 ;
        RECT -3.475 1.400 -3.305 2.350 ;
      LAYER mcon ;
        RECT -3.475 1.980 -3.305 2.150 ;
        RECT -3.475 1.620 -3.305 1.790 ;
      LAYER met1 ;
        RECT -3.520 1.395 -3.200 2.355 ;
      LAYER via ;
        RECT -3.490 1.915 -3.230 2.175 ;
        RECT -3.490 1.595 -3.230 1.855 ;
      LAYER met2 ;
        RECT -14.330 5.570 -12.515 7.350 ;
        RECT -13.135 1.025 -12.760 5.570 ;
        RECT -3.520 1.360 -3.200 2.355 ;
        RECT -3.725 1.165 -3.200 1.360 ;
        RECT -3.725 1.025 -3.315 1.165 ;
        RECT -13.135 0.765 -3.520 1.025 ;
    END
  END p100_SL
  PIN RE_BR0
    ANTENNADIFFAREA 4.200000 ;
    PORT
      LAYER li1 ;
        RECT 18.825 -2.820 18.995 2.530 ;
        RECT 18.725 -19.420 18.895 -14.070 ;
      LAYER mcon ;
        RECT 18.825 2.145 18.995 2.315 ;
        RECT 18.825 1.785 18.995 1.955 ;
        RECT 18.825 1.425 18.995 1.595 ;
        RECT 18.825 1.065 18.995 1.235 ;
        RECT 18.825 0.705 18.995 0.875 ;
        RECT 18.825 0.345 18.995 0.515 ;
        RECT 18.825 -0.015 18.995 0.155 ;
        RECT 18.825 -0.375 18.995 -0.205 ;
        RECT 18.825 -0.735 18.995 -0.565 ;
        RECT 18.825 -1.095 18.995 -0.925 ;
        RECT 18.825 -1.455 18.995 -1.285 ;
        RECT 18.825 -1.815 18.995 -1.645 ;
        RECT 18.825 -2.175 18.995 -2.005 ;
        RECT 18.825 -2.535 18.995 -2.365 ;
        RECT 18.725 -14.455 18.895 -14.285 ;
        RECT 18.725 -14.815 18.895 -14.645 ;
        RECT 18.725 -15.175 18.895 -15.005 ;
        RECT 18.725 -15.535 18.895 -15.365 ;
        RECT 18.725 -15.895 18.895 -15.725 ;
        RECT 18.725 -16.255 18.895 -16.085 ;
        RECT 18.725 -16.615 18.895 -16.445 ;
        RECT 18.725 -16.975 18.895 -16.805 ;
        RECT 18.725 -17.335 18.895 -17.165 ;
        RECT 18.725 -17.695 18.895 -17.525 ;
        RECT 18.725 -18.055 18.895 -17.885 ;
        RECT 18.725 -18.415 18.895 -18.245 ;
        RECT 18.725 -18.775 18.895 -18.605 ;
        RECT 18.725 -19.135 18.895 -18.965 ;
      LAYER met1 ;
        RECT 18.780 -3.080 19.100 2.535 ;
        RECT 18.780 -3.285 21.695 -3.080 ;
        RECT 21.415 -4.970 21.695 -3.285 ;
        RECT 18.680 -19.680 19.000 -14.065 ;
        RECT 18.680 -19.885 21.595 -19.680 ;
        RECT 21.315 -21.570 21.595 -19.885 ;
      LAYER via ;
        RECT 18.810 2.070 19.070 2.330 ;
        RECT 18.810 1.750 19.070 2.010 ;
        RECT 18.810 1.430 19.070 1.690 ;
        RECT 18.810 1.110 19.070 1.370 ;
        RECT 18.810 0.790 19.070 1.050 ;
        RECT 18.810 0.470 19.070 0.730 ;
        RECT 18.810 0.150 19.070 0.410 ;
        RECT 18.810 -0.170 19.070 0.090 ;
        RECT 18.810 -0.490 19.070 -0.230 ;
        RECT 18.810 -0.810 19.070 -0.550 ;
        RECT 18.810 -1.130 19.070 -0.870 ;
        RECT 18.810 -1.450 19.070 -1.190 ;
        RECT 18.810 -1.770 19.070 -1.510 ;
        RECT 18.810 -2.090 19.070 -1.830 ;
        RECT 18.810 -2.410 19.070 -2.150 ;
        RECT 18.810 -2.730 19.070 -2.470 ;
        RECT 21.420 -4.910 21.680 -4.650 ;
        RECT 18.710 -14.530 18.970 -14.270 ;
        RECT 18.710 -14.850 18.970 -14.590 ;
        RECT 18.710 -15.170 18.970 -14.910 ;
        RECT 18.710 -15.490 18.970 -15.230 ;
        RECT 18.710 -15.810 18.970 -15.550 ;
        RECT 18.710 -16.130 18.970 -15.870 ;
        RECT 18.710 -16.450 18.970 -16.190 ;
        RECT 18.710 -16.770 18.970 -16.510 ;
        RECT 18.710 -17.090 18.970 -16.830 ;
        RECT 18.710 -17.410 18.970 -17.150 ;
        RECT 18.710 -17.730 18.970 -17.470 ;
        RECT 18.710 -18.050 18.970 -17.790 ;
        RECT 18.710 -18.370 18.970 -18.110 ;
        RECT 18.710 -18.690 18.970 -18.430 ;
        RECT 18.710 -19.010 18.970 -18.750 ;
        RECT 18.710 -19.330 18.970 -19.070 ;
        RECT 21.320 -21.510 21.580 -21.250 ;
      LAYER met2 ;
        RECT 19.175 8.070 20.990 9.850 ;
        RECT 20.660 5.220 20.990 8.070 ;
        RECT 20.660 4.990 21.700 5.220 ;
        RECT 18.780 -2.815 19.100 2.535 ;
        RECT 21.195 -4.580 21.700 4.990 ;
        RECT 18.680 -19.415 19.000 -14.065 ;
        RECT 21.190 -14.970 21.695 -4.580 ;
        RECT 21.185 -16.000 21.695 -14.970 ;
        RECT 21.190 -21.180 21.695 -16.000 ;
        RECT 21.090 -21.570 21.695 -21.180 ;
    END
  END RE_BR0
  PIN BL0
    ANTENNADIFFAREA 0.244800 ;
    PORT
      LAYER li1 ;
        RECT 16.165 0.530 17.505 0.780 ;
        RECT 16.065 -16.070 17.405 -15.820 ;
      LAYER mcon ;
        RECT 16.475 0.570 16.645 0.740 ;
        RECT 16.375 -16.030 16.545 -15.860 ;
      LAYER met1 ;
        RECT 15.855 2.845 16.695 3.405 ;
        RECT 16.435 0.780 16.695 2.845 ;
        RECT 16.415 0.510 16.705 0.780 ;
        RECT 12.885 -4.200 13.160 -3.980 ;
        RECT 16.435 -4.200 16.695 0.510 ;
        RECT 12.885 -4.405 16.695 -4.200 ;
        RECT 15.755 -13.755 16.595 -13.195 ;
        RECT 16.335 -15.820 16.595 -13.755 ;
        RECT 16.315 -16.090 16.605 -15.820 ;
        RECT 12.785 -20.800 13.060 -20.580 ;
        RECT 16.335 -20.800 16.595 -16.090 ;
        RECT 12.785 -21.005 16.595 -20.800 ;
      LAYER via ;
        RECT 16.015 3.000 16.275 3.260 ;
        RECT 12.890 -4.350 13.150 -4.090 ;
        RECT 15.915 -13.600 16.175 -13.340 ;
        RECT 12.790 -20.950 13.050 -20.690 ;
      LAYER met2 ;
        RECT 11.355 8.070 13.170 9.850 ;
        RECT 12.880 -20.575 13.170 8.070 ;
        RECT 15.855 3.400 16.425 3.410 ;
        RECT 15.030 3.120 16.425 3.400 ;
        RECT 15.855 2.835 16.425 3.120 ;
        RECT 15.755 -13.200 16.325 -13.190 ;
        RECT 14.930 -13.480 16.325 -13.200 ;
        RECT 15.755 -13.765 16.325 -13.480 ;
        RECT 12.780 -21.000 13.170 -20.575 ;
    END
  END BL0
  PIN RE_BL0
    ANTENNADIFFAREA 4.200000 ;
    PORT
      LAYER li1 ;
        RECT 14.550 -2.820 14.720 2.530 ;
        RECT 14.450 -19.420 14.620 -14.070 ;
      LAYER mcon ;
        RECT 14.550 2.145 14.720 2.315 ;
        RECT 14.550 1.785 14.720 1.955 ;
        RECT 14.550 1.425 14.720 1.595 ;
        RECT 14.550 1.065 14.720 1.235 ;
        RECT 14.550 0.705 14.720 0.875 ;
        RECT 14.550 0.345 14.720 0.515 ;
        RECT 14.550 -0.015 14.720 0.155 ;
        RECT 14.550 -0.375 14.720 -0.205 ;
        RECT 14.550 -0.735 14.720 -0.565 ;
        RECT 14.550 -1.095 14.720 -0.925 ;
        RECT 14.550 -1.455 14.720 -1.285 ;
        RECT 14.550 -1.815 14.720 -1.645 ;
        RECT 14.550 -2.175 14.720 -2.005 ;
        RECT 14.550 -2.535 14.720 -2.365 ;
        RECT 14.450 -14.455 14.620 -14.285 ;
        RECT 14.450 -14.815 14.620 -14.645 ;
        RECT 14.450 -15.175 14.620 -15.005 ;
        RECT 14.450 -15.535 14.620 -15.365 ;
        RECT 14.450 -15.895 14.620 -15.725 ;
        RECT 14.450 -16.255 14.620 -16.085 ;
        RECT 14.450 -16.615 14.620 -16.445 ;
        RECT 14.450 -16.975 14.620 -16.805 ;
        RECT 14.450 -17.335 14.620 -17.165 ;
        RECT 14.450 -17.695 14.620 -17.525 ;
        RECT 14.450 -18.055 14.620 -17.885 ;
        RECT 14.450 -18.415 14.620 -18.245 ;
        RECT 14.450 -18.775 14.620 -18.605 ;
        RECT 14.450 -19.135 14.620 -18.965 ;
      LAYER met1 ;
        RECT 14.505 -2.465 14.825 2.535 ;
        RECT 12.245 -2.780 14.825 -2.465 ;
        RECT 12.245 -4.925 12.610 -2.780 ;
        RECT 14.505 -2.820 14.825 -2.780 ;
        RECT 14.405 -19.065 14.725 -14.065 ;
        RECT 12.145 -19.380 14.725 -19.065 ;
        RECT 12.145 -21.525 12.510 -19.380 ;
        RECT 14.405 -19.420 14.725 -19.380 ;
      LAYER via ;
        RECT 14.535 2.070 14.795 2.330 ;
        RECT 14.535 1.750 14.795 2.010 ;
        RECT 14.535 1.430 14.795 1.690 ;
        RECT 14.535 1.110 14.795 1.370 ;
        RECT 14.535 0.790 14.795 1.050 ;
        RECT 14.535 0.470 14.795 0.730 ;
        RECT 14.535 0.150 14.795 0.410 ;
        RECT 14.535 -0.170 14.795 0.090 ;
        RECT 14.535 -0.490 14.795 -0.230 ;
        RECT 14.535 -0.810 14.795 -0.550 ;
        RECT 14.535 -1.130 14.795 -0.870 ;
        RECT 14.535 -1.450 14.795 -1.190 ;
        RECT 14.535 -1.770 14.795 -1.510 ;
        RECT 14.535 -2.090 14.795 -1.830 ;
        RECT 14.535 -2.410 14.795 -2.150 ;
        RECT 14.535 -2.730 14.795 -2.470 ;
        RECT 12.315 -4.910 12.575 -4.650 ;
        RECT 14.435 -14.530 14.695 -14.270 ;
        RECT 14.435 -14.850 14.695 -14.590 ;
        RECT 14.435 -15.170 14.695 -14.910 ;
        RECT 14.435 -15.490 14.695 -15.230 ;
        RECT 14.435 -15.810 14.695 -15.550 ;
        RECT 14.435 -16.130 14.695 -15.870 ;
        RECT 14.435 -16.450 14.695 -16.190 ;
        RECT 14.435 -16.770 14.695 -16.510 ;
        RECT 14.435 -17.090 14.695 -16.830 ;
        RECT 14.435 -17.410 14.695 -17.150 ;
        RECT 14.435 -17.730 14.695 -17.470 ;
        RECT 14.435 -18.050 14.695 -17.790 ;
        RECT 14.435 -18.370 14.695 -18.110 ;
        RECT 14.435 -18.690 14.695 -18.430 ;
        RECT 14.435 -19.010 14.695 -18.750 ;
        RECT 14.435 -19.330 14.695 -19.070 ;
        RECT 12.215 -21.510 12.475 -21.250 ;
      LAYER met2 ;
        RECT 9.400 8.070 11.215 9.850 ;
        RECT 10.900 5.220 11.215 8.070 ;
        RECT 10.900 4.865 12.740 5.220 ;
        RECT 12.235 -4.970 12.740 4.865 ;
        RECT 14.505 -2.815 14.825 2.535 ;
        RECT 12.235 -14.970 12.640 -4.970 ;
        RECT 12.235 -16.000 12.740 -14.970 ;
        RECT 12.235 -21.180 12.640 -16.000 ;
        RECT 14.405 -19.415 14.725 -14.065 ;
        RECT 12.135 -21.570 12.740 -21.180 ;
    END
  END RE_BL0
  PIN BR0
    ANTENNADIFFAREA 0.244800 ;
    PORT
      LAYER li1 ;
        RECT 16.165 -1.620 17.505 -1.370 ;
        RECT 16.065 -18.220 17.405 -17.970 ;
      LAYER mcon ;
        RECT 17.015 -1.580 17.185 -1.410 ;
        RECT 16.915 -18.180 17.085 -18.010 ;
      LAYER met1 ;
        RECT 16.955 2.840 17.845 3.420 ;
        RECT 16.955 0.780 17.245 2.840 ;
        RECT 16.965 -1.350 17.225 0.780 ;
        RECT 16.955 -1.620 17.245 -1.350 ;
        RECT 16.965 -4.200 17.225 -1.620 ;
        RECT 20.660 -4.200 20.935 -3.980 ;
        RECT 16.965 -4.405 20.935 -4.200 ;
        RECT 16.965 -4.410 17.225 -4.405 ;
        RECT 16.855 -13.760 17.745 -13.180 ;
        RECT 16.855 -15.820 17.145 -13.760 ;
        RECT 16.865 -17.950 17.125 -15.820 ;
        RECT 16.855 -18.220 17.145 -17.950 ;
        RECT 16.865 -20.800 17.125 -18.220 ;
        RECT 20.560 -20.800 20.835 -20.580 ;
        RECT 16.865 -21.005 20.835 -20.800 ;
        RECT 16.865 -21.010 17.125 -21.005 ;
      LAYER via ;
        RECT 17.425 2.990 17.685 3.250 ;
        RECT 20.665 -4.350 20.925 -4.090 ;
        RECT 17.325 -13.610 17.585 -13.350 ;
        RECT 20.565 -20.950 20.825 -20.690 ;
      LAYER met2 ;
        RECT 17.220 8.070 19.035 9.850 ;
        RECT 18.725 4.700 19.035 8.070 ;
        RECT 18.725 4.515 20.945 4.700 ;
        RECT 17.250 3.150 18.985 3.420 ;
        RECT 17.250 2.845 17.840 3.150 ;
        RECT 17.150 -13.450 18.885 -13.180 ;
        RECT 17.150 -13.755 17.740 -13.450 ;
        RECT 20.655 -20.575 20.945 4.515 ;
        RECT 20.555 -21.000 20.945 -20.575 ;
    END
  END BR0
  PIN p1T1R_TE
    PORT
      LAYER met2 ;
        RECT -8.465 5.570 -6.650 7.350 ;
        RECT -7.065 3.245 -6.650 5.570 ;
        RECT -7.065 3.240 -0.860 3.245 ;
        RECT -7.065 2.920 -4.530 3.240 ;
        RECT -4.210 2.920 -3.315 3.240 ;
        RECT -2.995 2.920 -2.260 3.240 ;
        RECT -1.940 2.920 -1.225 3.240 ;
        RECT -0.905 2.920 -0.860 3.240 ;
        RECT -7.065 2.900 -0.860 2.920 ;
    END
  END p1T1R_TE
  PIN p1R_SL
    PORT
      LAYER met1 ;
        RECT -5.710 4.435 -4.410 4.695 ;
      LAYER via ;
        RECT -5.670 4.435 -5.410 4.695 ;
      LAYER met2 ;
        RECT -6.510 5.570 -4.695 7.350 ;
        RECT -6.000 4.300 -5.055 5.570 ;
    END
  END p1R_SL
  PIN p1R_TE
    PORT
      LAYER met2 ;
        RECT -4.555 5.570 -2.740 7.350 ;
        RECT -4.555 4.725 -4.000 5.570 ;
        RECT -4.410 4.405 -4.000 4.725 ;
    END
  END p1R_TE
  PIN BR1
    ANTENNADIFFAREA 0.244800 ;
    PORT
      LAYER li1 ;
        RECT 36.415 -1.620 37.755 -1.370 ;
        RECT 36.315 -18.220 37.655 -17.970 ;
      LAYER mcon ;
        RECT 37.265 -1.580 37.435 -1.410 ;
        RECT 37.165 -18.180 37.335 -18.010 ;
      LAYER met1 ;
        RECT 37.205 2.840 38.095 3.420 ;
        RECT 37.205 0.780 37.495 2.840 ;
        RECT 37.215 -1.350 37.475 0.780 ;
        RECT 37.205 -1.620 37.495 -1.350 ;
        RECT 37.215 -4.200 37.475 -1.620 ;
        RECT 40.910 -4.200 41.185 -3.980 ;
        RECT 37.215 -4.405 41.185 -4.200 ;
        RECT 37.215 -4.410 37.475 -4.405 ;
        RECT 37.105 -13.760 37.995 -13.180 ;
        RECT 37.105 -15.820 37.395 -13.760 ;
        RECT 37.115 -17.950 37.375 -15.820 ;
        RECT 37.105 -18.220 37.395 -17.950 ;
        RECT 37.115 -20.800 37.375 -18.220 ;
        RECT 40.810 -20.800 41.085 -20.580 ;
        RECT 37.115 -21.005 41.085 -20.800 ;
        RECT 37.115 -21.010 37.375 -21.005 ;
      LAYER via ;
        RECT 37.675 2.990 37.935 3.250 ;
        RECT 40.915 -4.350 41.175 -4.090 ;
        RECT 37.575 -13.610 37.835 -13.350 ;
        RECT 40.815 -20.950 41.075 -20.690 ;
      LAYER met2 ;
        RECT 35.290 8.070 37.105 9.850 ;
        RECT 36.890 4.070 37.105 8.070 ;
        RECT 36.890 3.925 41.190 4.070 ;
        RECT 37.500 3.150 39.235 3.420 ;
        RECT 37.500 2.845 38.090 3.150 ;
        RECT 40.900 -3.975 41.190 3.925 ;
        RECT 37.400 -13.450 39.135 -13.180 ;
        RECT 37.400 -13.755 37.990 -13.450 ;
        RECT 40.905 -20.575 41.195 -3.975 ;
        RECT 40.805 -21.000 41.195 -20.575 ;
    END
  END BR1
  PIN RE_BR1
    ANTENNADIFFAREA 4.200000 ;
    PORT
      LAYER li1 ;
        RECT 39.075 -2.820 39.245 2.530 ;
        RECT 38.975 -19.420 39.145 -14.070 ;
      LAYER mcon ;
        RECT 39.075 2.145 39.245 2.315 ;
        RECT 39.075 1.785 39.245 1.955 ;
        RECT 39.075 1.425 39.245 1.595 ;
        RECT 39.075 1.065 39.245 1.235 ;
        RECT 39.075 0.705 39.245 0.875 ;
        RECT 39.075 0.345 39.245 0.515 ;
        RECT 39.075 -0.015 39.245 0.155 ;
        RECT 39.075 -0.375 39.245 -0.205 ;
        RECT 39.075 -0.735 39.245 -0.565 ;
        RECT 39.075 -1.095 39.245 -0.925 ;
        RECT 39.075 -1.455 39.245 -1.285 ;
        RECT 39.075 -1.815 39.245 -1.645 ;
        RECT 39.075 -2.175 39.245 -2.005 ;
        RECT 39.075 -2.535 39.245 -2.365 ;
        RECT 38.975 -14.455 39.145 -14.285 ;
        RECT 38.975 -14.815 39.145 -14.645 ;
        RECT 38.975 -15.175 39.145 -15.005 ;
        RECT 38.975 -15.535 39.145 -15.365 ;
        RECT 38.975 -15.895 39.145 -15.725 ;
        RECT 38.975 -16.255 39.145 -16.085 ;
        RECT 38.975 -16.615 39.145 -16.445 ;
        RECT 38.975 -16.975 39.145 -16.805 ;
        RECT 38.975 -17.335 39.145 -17.165 ;
        RECT 38.975 -17.695 39.145 -17.525 ;
        RECT 38.975 -18.055 39.145 -17.885 ;
        RECT 38.975 -18.415 39.145 -18.245 ;
        RECT 38.975 -18.775 39.145 -18.605 ;
        RECT 38.975 -19.135 39.145 -18.965 ;
      LAYER met1 ;
        RECT 39.030 -3.080 39.350 2.535 ;
        RECT 39.030 -3.285 41.945 -3.080 ;
        RECT 41.665 -4.970 41.945 -3.285 ;
        RECT 38.930 -19.680 39.250 -14.065 ;
        RECT 38.930 -19.885 41.845 -19.680 ;
        RECT 41.565 -21.570 41.845 -19.885 ;
      LAYER via ;
        RECT 39.060 2.070 39.320 2.330 ;
        RECT 39.060 1.750 39.320 2.010 ;
        RECT 39.060 1.430 39.320 1.690 ;
        RECT 39.060 1.110 39.320 1.370 ;
        RECT 39.060 0.790 39.320 1.050 ;
        RECT 39.060 0.470 39.320 0.730 ;
        RECT 39.060 0.150 39.320 0.410 ;
        RECT 39.060 -0.170 39.320 0.090 ;
        RECT 39.060 -0.490 39.320 -0.230 ;
        RECT 39.060 -0.810 39.320 -0.550 ;
        RECT 39.060 -1.130 39.320 -0.870 ;
        RECT 39.060 -1.450 39.320 -1.190 ;
        RECT 39.060 -1.770 39.320 -1.510 ;
        RECT 39.060 -2.090 39.320 -1.830 ;
        RECT 39.060 -2.410 39.320 -2.150 ;
        RECT 39.060 -2.730 39.320 -2.470 ;
        RECT 41.670 -4.910 41.930 -4.650 ;
        RECT 38.960 -14.530 39.220 -14.270 ;
        RECT 38.960 -14.850 39.220 -14.590 ;
        RECT 38.960 -15.170 39.220 -14.910 ;
        RECT 38.960 -15.490 39.220 -15.230 ;
        RECT 38.960 -15.810 39.220 -15.550 ;
        RECT 38.960 -16.130 39.220 -15.870 ;
        RECT 38.960 -16.450 39.220 -16.190 ;
        RECT 38.960 -16.770 39.220 -16.510 ;
        RECT 38.960 -17.090 39.220 -16.830 ;
        RECT 38.960 -17.410 39.220 -17.150 ;
        RECT 38.960 -17.730 39.220 -17.470 ;
        RECT 38.960 -18.050 39.220 -17.790 ;
        RECT 38.960 -18.370 39.220 -18.110 ;
        RECT 38.960 -18.690 39.220 -18.430 ;
        RECT 38.960 -19.010 39.220 -18.750 ;
        RECT 38.960 -19.330 39.220 -19.070 ;
        RECT 41.570 -21.510 41.830 -21.250 ;
      LAYER met2 ;
        RECT 37.245 8.070 39.060 9.850 ;
        RECT 38.795 4.395 39.060 8.070 ;
        RECT 38.795 4.210 41.945 4.395 ;
        RECT 39.030 -2.815 39.350 2.535 ;
        RECT 38.930 -19.415 39.250 -14.065 ;
        RECT 41.440 -14.970 41.945 4.210 ;
        RECT 41.435 -16.000 41.945 -14.970 ;
        RECT 41.440 -21.180 41.945 -16.000 ;
        RECT 41.340 -21.570 41.945 -21.180 ;
    END
  END RE_BR1
  PIN BL1
    ANTENNADIFFAREA 0.244800 ;
    PORT
      LAYER li1 ;
        RECT 36.415 0.530 37.755 0.780 ;
        RECT 36.315 -16.070 37.655 -15.820 ;
      LAYER mcon ;
        RECT 36.725 0.570 36.895 0.740 ;
        RECT 36.625 -16.030 36.795 -15.860 ;
      LAYER met1 ;
        RECT 36.105 2.845 36.945 3.405 ;
        RECT 36.685 0.780 36.945 2.845 ;
        RECT 36.665 0.510 36.955 0.780 ;
        RECT 33.135 -4.200 33.410 -3.980 ;
        RECT 36.685 -4.200 36.945 0.510 ;
        RECT 33.135 -4.405 36.945 -4.200 ;
        RECT 36.005 -13.755 36.845 -13.195 ;
        RECT 36.585 -15.820 36.845 -13.755 ;
        RECT 36.565 -16.090 36.855 -15.820 ;
        RECT 33.035 -20.800 33.310 -20.580 ;
        RECT 36.585 -20.800 36.845 -16.090 ;
        RECT 33.035 -21.005 36.845 -20.800 ;
      LAYER via ;
        RECT 36.265 3.000 36.525 3.260 ;
        RECT 33.140 -4.350 33.400 -4.090 ;
        RECT 36.165 -13.600 36.425 -13.340 ;
        RECT 33.040 -20.950 33.300 -20.690 ;
      LAYER met2 ;
        RECT 33.335 8.070 35.150 9.850 ;
        RECT 33.335 5.220 33.735 8.070 ;
        RECT 33.125 5.055 33.735 5.220 ;
        RECT 33.125 -3.975 33.415 5.055 ;
        RECT 36.105 3.400 36.675 3.410 ;
        RECT 35.280 3.120 36.675 3.400 ;
        RECT 36.105 2.835 36.675 3.120 ;
        RECT 33.130 -20.575 33.420 -3.975 ;
        RECT 36.005 -13.200 36.575 -13.190 ;
        RECT 35.180 -13.480 36.575 -13.200 ;
        RECT 36.005 -13.765 36.575 -13.480 ;
        RECT 33.030 -21.000 33.420 -20.575 ;
    END
  END BL1
  PIN RE_BL1
    ANTENNADIFFAREA 4.200000 ;
    PORT
      LAYER li1 ;
        RECT 34.800 -2.820 34.970 2.530 ;
        RECT 34.700 -19.420 34.870 -14.070 ;
      LAYER mcon ;
        RECT 34.800 2.145 34.970 2.315 ;
        RECT 34.800 1.785 34.970 1.955 ;
        RECT 34.800 1.425 34.970 1.595 ;
        RECT 34.800 1.065 34.970 1.235 ;
        RECT 34.800 0.705 34.970 0.875 ;
        RECT 34.800 0.345 34.970 0.515 ;
        RECT 34.800 -0.015 34.970 0.155 ;
        RECT 34.800 -0.375 34.970 -0.205 ;
        RECT 34.800 -0.735 34.970 -0.565 ;
        RECT 34.800 -1.095 34.970 -0.925 ;
        RECT 34.800 -1.455 34.970 -1.285 ;
        RECT 34.800 -1.815 34.970 -1.645 ;
        RECT 34.800 -2.175 34.970 -2.005 ;
        RECT 34.800 -2.535 34.970 -2.365 ;
        RECT 34.700 -14.455 34.870 -14.285 ;
        RECT 34.700 -14.815 34.870 -14.645 ;
        RECT 34.700 -15.175 34.870 -15.005 ;
        RECT 34.700 -15.535 34.870 -15.365 ;
        RECT 34.700 -15.895 34.870 -15.725 ;
        RECT 34.700 -16.255 34.870 -16.085 ;
        RECT 34.700 -16.615 34.870 -16.445 ;
        RECT 34.700 -16.975 34.870 -16.805 ;
        RECT 34.700 -17.335 34.870 -17.165 ;
        RECT 34.700 -17.695 34.870 -17.525 ;
        RECT 34.700 -18.055 34.870 -17.885 ;
        RECT 34.700 -18.415 34.870 -18.245 ;
        RECT 34.700 -18.775 34.870 -18.605 ;
        RECT 34.700 -19.135 34.870 -18.965 ;
      LAYER met1 ;
        RECT 34.755 -2.465 35.075 2.535 ;
        RECT 32.495 -2.780 35.075 -2.465 ;
        RECT 32.495 -4.925 32.860 -2.780 ;
        RECT 34.755 -2.820 35.075 -2.780 ;
        RECT 34.655 -19.065 34.975 -14.065 ;
        RECT 32.395 -19.380 34.975 -19.065 ;
        RECT 32.395 -21.525 32.760 -19.380 ;
        RECT 34.655 -19.420 34.975 -19.380 ;
      LAYER via ;
        RECT 34.785 2.070 35.045 2.330 ;
        RECT 34.785 1.750 35.045 2.010 ;
        RECT 34.785 1.430 35.045 1.690 ;
        RECT 34.785 1.110 35.045 1.370 ;
        RECT 34.785 0.790 35.045 1.050 ;
        RECT 34.785 0.470 35.045 0.730 ;
        RECT 34.785 0.150 35.045 0.410 ;
        RECT 34.785 -0.170 35.045 0.090 ;
        RECT 34.785 -0.490 35.045 -0.230 ;
        RECT 34.785 -0.810 35.045 -0.550 ;
        RECT 34.785 -1.130 35.045 -0.870 ;
        RECT 34.785 -1.450 35.045 -1.190 ;
        RECT 34.785 -1.770 35.045 -1.510 ;
        RECT 34.785 -2.090 35.045 -1.830 ;
        RECT 34.785 -2.410 35.045 -2.150 ;
        RECT 34.785 -2.730 35.045 -2.470 ;
        RECT 32.565 -4.910 32.825 -4.650 ;
        RECT 34.685 -14.530 34.945 -14.270 ;
        RECT 34.685 -14.850 34.945 -14.590 ;
        RECT 34.685 -15.170 34.945 -14.910 ;
        RECT 34.685 -15.490 34.945 -15.230 ;
        RECT 34.685 -15.810 34.945 -15.550 ;
        RECT 34.685 -16.130 34.945 -15.870 ;
        RECT 34.685 -16.450 34.945 -16.190 ;
        RECT 34.685 -16.770 34.945 -16.510 ;
        RECT 34.685 -17.090 34.945 -16.830 ;
        RECT 34.685 -17.410 34.945 -17.150 ;
        RECT 34.685 -17.730 34.945 -17.470 ;
        RECT 34.685 -18.050 34.945 -17.790 ;
        RECT 34.685 -18.370 34.945 -18.110 ;
        RECT 34.685 -18.690 34.945 -18.430 ;
        RECT 34.685 -19.010 34.945 -18.750 ;
        RECT 34.685 -19.330 34.945 -19.070 ;
        RECT 32.465 -21.510 32.725 -21.250 ;
      LAYER met2 ;
        RECT 31.180 8.070 32.995 9.850 ;
        RECT 32.480 -4.580 32.985 8.070 ;
        RECT 34.755 -2.815 35.075 2.535 ;
        RECT 32.485 -4.970 32.990 -4.580 ;
        RECT 32.485 -14.970 32.890 -4.970 ;
        RECT 32.485 -16.000 32.990 -14.970 ;
        RECT 32.485 -21.180 32.890 -16.000 ;
        RECT 34.655 -19.415 34.975 -14.065 ;
        RECT 32.385 -21.570 32.990 -21.180 ;
    END
  END RE_BL1
  PIN RE_WL1
    ANTENNAGATEAREA 4.200000 ;
    PORT
      LAYER li1 ;
        RECT 45.380 -20.675 45.780 -20.385 ;
        RECT 10.750 -20.845 22.820 -20.675 ;
        RECT 31.000 -20.845 45.780 -20.675 ;
        RECT 14.630 -21.525 14.985 -20.845 ;
        RECT 18.905 -21.525 19.260 -20.845 ;
        RECT 34.880 -21.525 35.235 -20.845 ;
        RECT 39.155 -21.525 39.510 -20.845 ;
      LAYER mcon ;
        RECT 22.565 -20.845 22.735 -20.675 ;
        RECT 31.110 -20.845 31.280 -20.675 ;
        RECT 45.485 -20.680 45.655 -20.510 ;
      LAYER met1 ;
        RECT 22.455 -20.995 31.365 -20.630 ;
        RECT 45.380 -20.805 45.780 -20.385 ;
      LAYER via ;
        RECT 45.455 -20.720 45.715 -20.460 ;
      LAYER met2 ;
        RECT 45.065 8.070 46.880 9.850 ;
        RECT 45.380 -20.845 45.780 8.070 ;
    END
  END RE_WL1
  PIN RE_WL0
    ANTENNAGATEAREA 4.200000 ;
    PORT
      LAYER li1 ;
        RECT 42.970 -4.075 43.370 -3.825 ;
        RECT 10.850 -4.245 22.725 -4.075 ;
        RECT 31.100 -4.245 45.870 -4.075 ;
        RECT 14.730 -4.925 15.085 -4.245 ;
        RECT 19.005 -4.925 19.360 -4.245 ;
        RECT 34.980 -4.925 35.335 -4.245 ;
        RECT 39.255 -4.925 39.610 -4.245 ;
      LAYER mcon ;
        RECT 22.470 -4.245 22.640 -4.075 ;
        RECT 31.210 -4.245 31.380 -4.075 ;
        RECT 43.075 -4.120 43.245 -3.950 ;
      LAYER met1 ;
        RECT 22.360 -4.395 31.465 -4.030 ;
        RECT 42.970 -4.245 43.370 -3.825 ;
      LAYER via ;
        RECT 43.045 -4.160 43.305 -3.900 ;
      LAYER met2 ;
        RECT 41.155 8.070 42.970 9.850 ;
        RECT 42.590 5.270 42.970 8.070 ;
        RECT 42.590 4.910 43.370 5.270 ;
        RECT 42.970 -4.245 43.370 4.910 ;
    END
  END RE_WL0
  PIN WL1
    ANTENNAGATEAREA 0.216000 ;
    PORT
      LAYER li1 ;
        RECT 15.290 -20.215 15.605 -19.660 ;
        RECT 35.540 -20.215 35.855 -19.660 ;
        RECT 43.820 -20.215 44.220 -19.925 ;
        RECT 10.750 -20.385 22.820 -20.215 ;
        RECT 31.000 -20.385 44.220 -20.215 ;
      LAYER mcon ;
        RECT 22.565 -20.385 22.735 -20.215 ;
        RECT 31.110 -20.385 31.280 -20.215 ;
        RECT 43.925 -20.220 44.095 -20.050 ;
      LAYER met1 ;
        RECT 22.455 -20.430 31.365 -20.040 ;
        RECT 43.820 -20.345 44.220 -19.925 ;
      LAYER via ;
        RECT 43.895 -20.260 44.155 -20.000 ;
      LAYER met2 ;
        RECT 43.110 8.070 44.925 9.850 ;
        RECT 43.820 -20.385 44.220 8.070 ;
    END
  END WL1
  PIN WL0
    ANTENNAGATEAREA 0.216000 ;
    PORT
      LAYER li1 ;
        RECT 15.390 -3.615 15.705 -3.060 ;
        RECT 35.640 -3.615 35.955 -3.060 ;
        RECT 42.270 -3.615 42.670 -3.365 ;
        RECT 10.850 -3.785 22.725 -3.615 ;
        RECT 31.100 -3.785 42.670 -3.615 ;
      LAYER mcon ;
        RECT 22.470 -3.785 22.640 -3.615 ;
        RECT 31.210 -3.785 31.380 -3.615 ;
        RECT 42.375 -3.660 42.545 -3.490 ;
      LAYER met1 ;
        RECT 22.360 -3.830 31.465 -3.440 ;
        RECT 42.270 -3.785 42.670 -3.365 ;
      LAYER via ;
        RECT 42.345 -3.700 42.605 -3.440 ;
      LAYER met2 ;
        RECT 39.200 8.070 41.015 9.850 ;
        RECT 40.605 4.695 41.010 8.070 ;
        RECT 40.605 4.535 42.670 4.695 ;
        RECT 42.270 -3.785 42.670 4.535 ;
    END
  END WL0
  PIN pVDD_HEADER0
    ANTENNAGATEAREA 0.108000 ;
    PORT
      LAYER li1 ;
        RECT 15.865 5.500 16.425 5.785 ;
        RECT 36.115 5.500 36.675 5.785 ;
      LAYER mcon ;
        RECT 16.200 5.565 16.370 5.735 ;
        RECT 36.450 5.565 36.620 5.735 ;
      LAYER met1 ;
        RECT 15.825 5.465 36.755 5.935 ;
      LAYER via ;
        RECT 23.375 5.555 23.635 5.815 ;
      LAYER met2 ;
        RECT 22.730 8.070 24.545 9.850 ;
        RECT 23.225 5.365 23.790 8.070 ;
    END
  END pVDD_HEADER0
  PIN pGND_HEADER0
    ANTENNAGATEAREA 0.108000 ;
    PORT
      LAYER li1 ;
        RECT 17.460 4.875 18.020 5.160 ;
        RECT 37.710 4.875 38.270 5.160 ;
      LAYER mcon ;
        RECT 17.795 4.940 17.965 5.110 ;
        RECT 38.045 4.940 38.215 5.110 ;
      LAYER met1 ;
        RECT 17.380 4.825 31.560 5.225 ;
        RECT 37.945 5.160 38.280 6.650 ;
        RECT 37.910 4.875 38.345 5.160 ;
      LAYER via ;
        RECT 37.985 6.355 38.245 6.615 ;
        RECT 25.500 4.885 25.760 5.145 ;
        RECT 31.180 4.900 31.440 5.160 ;
      LAYER met2 ;
        RECT 24.685 8.070 26.500 9.850 ;
        RECT 25.345 4.090 25.910 8.070 ;
        RECT 31.100 4.830 31.965 6.795 ;
        RECT 37.635 6.120 38.365 6.890 ;
      LAYER via2 ;
        RECT 31.370 6.385 31.650 6.665 ;
        RECT 37.970 6.345 38.250 6.625 ;
      LAYER met3 ;
        RECT 31.100 6.180 38.335 6.795 ;
    END
  END pGND_HEADER0
  PIN pVDD_HEADER1
    ANTENNAGATEAREA 0.108000 ;
    PORT
      LAYER li1 ;
        RECT 15.765 -11.100 16.325 -10.815 ;
        RECT 36.015 -11.100 36.575 -10.815 ;
      LAYER mcon ;
        RECT 16.100 -11.035 16.270 -10.865 ;
        RECT 36.350 -11.035 36.520 -10.865 ;
      LAYER met1 ;
        RECT 15.725 -10.815 36.425 -10.685 ;
        RECT 15.725 -11.100 36.650 -10.815 ;
        RECT 15.725 -11.155 36.425 -11.100 ;
      LAYER via ;
        RECT 27.775 -11.065 28.035 -10.805 ;
      LAYER met2 ;
        RECT 26.640 8.070 28.455 9.850 ;
        RECT 27.625 -11.255 28.190 8.070 ;
    END
  END pVDD_HEADER1
  PIN pGND_HEADER1
    ANTENNAGATEAREA 0.108000 ;
    PORT
      LAYER li1 ;
        RECT 17.360 -11.725 17.920 -11.440 ;
        RECT 37.610 -11.725 38.170 -11.440 ;
      LAYER mcon ;
        RECT 17.695 -11.660 17.865 -11.490 ;
        RECT 37.945 -11.660 38.115 -11.490 ;
      LAYER met1 ;
        RECT 37.710 -10.425 38.555 -9.660 ;
        RECT 17.280 -11.775 30.110 -11.375 ;
        RECT 37.810 -11.725 38.245 -10.425 ;
      LAYER via ;
        RECT 38.000 -10.175 38.260 -9.915 ;
        RECT 29.690 -11.700 29.950 -11.440 ;
      LAYER met2 ;
        RECT 28.595 8.070 30.410 9.850 ;
        RECT 29.545 -12.510 30.110 8.070 ;
        RECT 37.710 -10.425 38.555 -9.660 ;
      LAYER via2 ;
        RECT 29.685 -10.185 29.965 -9.905 ;
        RECT 37.985 -10.185 38.265 -9.905 ;
      LAYER met3 ;
        RECT 29.545 -10.250 38.435 -9.850 ;
    END
  END pGND_HEADER1
  PIN vssd1
    ANTENNADIFFAREA 0.432000 ;
    PORT
      LAYER li1 ;
        RECT 17.290 4.315 17.460 4.645 ;
        RECT 37.540 4.315 37.710 4.645 ;
        RECT -6.145 3.565 -2.240 4.025 ;
        RECT -6.145 -1.395 -5.315 3.565 ;
        RECT -6.145 -2.230 -2.155 -1.395 ;
        RECT 17.490 -2.505 17.750 -1.925 ;
        RECT 37.740 -2.505 38.000 -1.925 ;
        RECT 17.190 -12.285 17.360 -11.955 ;
        RECT 37.440 -12.285 37.610 -11.955 ;
        RECT 17.390 -19.105 17.650 -18.525 ;
        RECT 37.640 -19.105 37.900 -18.525 ;
      LAYER mcon ;
        RECT 17.290 4.395 17.460 4.565 ;
        RECT 37.540 4.395 37.710 4.565 ;
        RECT -5.460 3.720 -5.290 3.890 ;
        RECT -4.990 3.715 -4.820 3.885 ;
        RECT -4.465 3.705 -4.295 3.875 ;
        RECT -3.995 3.700 -3.825 3.870 ;
        RECT -3.570 3.710 -3.400 3.880 ;
        RECT -3.100 3.705 -2.930 3.875 ;
        RECT -2.575 3.695 -2.405 3.865 ;
        RECT -5.840 3.390 -5.670 3.560 ;
        RECT -5.840 2.920 -5.670 3.090 ;
        RECT -5.850 2.385 -5.680 2.555 ;
        RECT -5.845 1.870 -5.675 2.040 ;
        RECT -5.845 1.130 -5.675 1.300 ;
        RECT -5.835 0.590 -5.665 0.760 ;
        RECT -5.845 -0.005 -5.675 0.165 ;
        RECT -5.845 -0.570 -5.675 -0.400 ;
        RECT -5.825 -1.230 -5.655 -1.060 ;
        RECT -5.835 -1.825 -5.665 -1.655 ;
        RECT -5.365 -1.830 -5.195 -1.660 ;
        RECT -4.840 -1.840 -4.670 -1.670 ;
        RECT -4.370 -1.845 -4.200 -1.675 ;
        RECT -3.945 -1.835 -3.775 -1.665 ;
        RECT -3.475 -1.840 -3.305 -1.670 ;
        RECT -2.950 -1.850 -2.780 -1.680 ;
        RECT 17.540 -2.360 17.710 -2.190 ;
        RECT 37.790 -2.360 37.960 -2.190 ;
        RECT 17.190 -12.205 17.360 -12.035 ;
        RECT 37.440 -12.205 37.610 -12.035 ;
        RECT 17.440 -18.960 17.610 -18.790 ;
        RECT 37.690 -18.960 37.860 -18.790 ;
      LAYER met1 ;
        RECT 17.060 14.305 18.880 15.100 ;
        RECT 8.170 14.085 18.880 14.305 ;
        RECT 8.170 6.285 8.425 14.085 ;
        RECT 17.060 13.320 18.880 14.085 ;
        RECT -2.605 6.060 8.425 6.285 ;
        RECT -2.605 3.965 -2.330 6.060 ;
        RECT 17.215 4.310 17.565 4.645 ;
        RECT 37.465 4.310 37.815 4.645 ;
        RECT -5.950 3.625 -2.330 3.965 ;
        RECT -5.950 -1.595 -5.560 3.625 ;
        RECT -5.950 -1.960 -2.355 -1.595 ;
        RECT 17.485 -3.855 17.745 -2.005 ;
        RECT 20.020 -3.855 20.380 -3.685 ;
        RECT 17.485 -4.060 20.380 -3.855 ;
        RECT 37.735 -3.855 37.995 -2.005 ;
        RECT 40.270 -3.855 40.630 -3.685 ;
        RECT 37.735 -4.060 40.630 -3.855 ;
        RECT 20.020 -9.500 40.635 -9.130 ;
        RECT 17.115 -12.290 17.465 -11.955 ;
        RECT 37.365 -12.290 37.715 -11.955 ;
        RECT 17.385 -20.455 17.645 -18.605 ;
        RECT 19.920 -20.455 20.280 -20.285 ;
        RECT 17.385 -20.660 20.280 -20.455 ;
        RECT 37.635 -20.455 37.895 -18.605 ;
        RECT 40.170 -20.455 40.530 -20.285 ;
        RECT 37.635 -20.660 40.530 -20.455 ;
      LAYER via ;
        RECT 17.330 14.380 17.590 14.640 ;
        RECT 17.855 14.405 18.115 14.665 ;
        RECT 18.375 14.405 18.635 14.665 ;
        RECT 17.330 14.060 17.590 14.320 ;
        RECT 17.855 14.085 18.115 14.345 ;
        RECT 18.375 14.085 18.635 14.345 ;
        RECT 17.330 13.740 17.590 14.000 ;
        RECT 17.855 13.765 18.115 14.025 ;
        RECT 18.375 13.765 18.635 14.025 ;
        RECT 17.265 4.335 17.525 4.595 ;
        RECT 37.525 4.350 37.785 4.610 ;
        RECT 20.065 -3.995 20.325 -3.735 ;
        RECT 40.315 -3.995 40.575 -3.735 ;
        RECT 20.065 -9.435 20.325 -9.175 ;
        RECT 40.320 -9.440 40.580 -9.180 ;
        RECT 17.140 -12.255 17.400 -11.995 ;
        RECT 37.405 -12.250 37.665 -11.990 ;
        RECT 19.965 -20.595 20.225 -20.335 ;
        RECT 40.215 -20.595 40.475 -20.335 ;
      LAYER met2 ;
        RECT 16.750 13.320 18.900 15.100 ;
        RECT 16.750 4.015 17.080 13.320 ;
        RECT 17.225 4.250 17.720 4.930 ;
        RECT 37.435 4.275 37.890 4.700 ;
        RECT 16.750 3.670 20.385 4.015 ;
        RECT 16.925 -12.500 17.500 -11.820 ;
        RECT 20.020 -20.280 20.385 3.670 ;
        RECT 40.265 -3.680 40.630 3.570 ;
        RECT 37.145 -12.700 37.885 -11.735 ;
        RECT 40.270 -20.280 40.635 -3.680 ;
        RECT 19.920 -20.660 20.385 -20.280 ;
        RECT 40.170 -20.660 40.635 -20.280 ;
      LAYER via2 ;
        RECT 17.140 14.345 17.420 14.625 ;
        RECT 17.625 14.345 17.905 14.625 ;
        RECT 18.135 14.345 18.415 14.625 ;
        RECT 17.140 13.930 17.420 14.210 ;
        RECT 17.625 13.930 17.905 14.210 ;
        RECT 18.135 13.930 18.415 14.210 ;
        RECT 17.140 13.490 17.420 13.770 ;
        RECT 17.625 13.490 17.905 13.770 ;
        RECT 18.135 13.490 18.415 13.770 ;
        RECT 17.255 4.325 17.535 4.605 ;
        RECT 37.520 4.325 37.800 4.605 ;
        RECT 16.955 -12.425 17.235 -12.145 ;
        RECT 37.395 -12.260 37.675 -11.980 ;
      LAYER met3 ;
        RECT 16.855 13.320 18.675 15.100 ;
        RECT 17.225 4.250 37.905 4.665 ;
        RECT 16.925 -12.345 17.420 -11.820 ;
        RECT 37.370 -12.345 37.700 -11.920 ;
        RECT 16.925 -12.825 37.700 -12.345 ;
        RECT 17.420 -12.830 37.700 -12.825 ;
      LAYER via3 ;
        RECT 17.120 14.325 17.440 14.645 ;
        RECT 17.605 14.325 17.925 14.645 ;
        RECT 18.115 14.325 18.435 14.645 ;
        RECT 17.120 13.910 17.440 14.230 ;
        RECT 17.605 13.910 17.925 14.230 ;
        RECT 18.115 13.910 18.435 14.230 ;
        RECT 17.120 13.470 17.440 13.790 ;
        RECT 17.605 13.470 17.925 13.790 ;
        RECT 18.115 13.470 18.435 13.790 ;
        RECT 17.235 4.305 17.555 4.625 ;
        RECT 16.935 -12.445 17.255 -12.125 ;
      LAYER met4 ;
        RECT 16.910 -72.000 18.650 165.250 ;
    END
  END vssd1
  PIN vccd1
    ANTENNADIFFAREA 1.132100 ;
    PORT
      LAYER nwell ;
        RECT 15.530 5.470 16.530 5.830 ;
        RECT 35.780 5.470 36.780 5.830 ;
        RECT 14.860 4.440 16.530 5.470 ;
        RECT 34.910 4.370 36.780 5.470 ;
        RECT 15.715 -2.505 16.695 0.780 ;
        RECT 35.965 -2.505 36.945 0.780 ;
        RECT 15.430 -11.130 16.430 -10.770 ;
        RECT 35.680 -11.130 36.680 -10.770 ;
        RECT 14.715 -12.075 16.430 -11.130 ;
        RECT 34.885 -12.245 36.680 -11.130 ;
        RECT 15.615 -19.105 16.595 -15.820 ;
        RECT 35.865 -19.105 36.845 -15.820 ;
      LAYER li1 ;
        RECT 14.950 4.940 15.865 5.270 ;
        RECT 35.265 4.940 36.115 5.270 ;
        RECT 15.915 -2.505 16.175 -1.925 ;
        RECT 36.165 -2.505 36.425 -1.925 ;
        RECT 14.840 -11.660 15.765 -11.330 ;
        RECT 35.010 -11.660 36.015 -11.330 ;
        RECT 15.815 -19.105 16.075 -18.525 ;
        RECT 36.065 -19.105 36.325 -18.525 ;
      LAYER mcon ;
        RECT 15.695 5.020 15.865 5.190 ;
        RECT 35.945 5.020 36.115 5.190 ;
        RECT 15.965 -2.360 16.135 -2.190 ;
        RECT 36.215 -2.360 36.385 -2.190 ;
        RECT 15.595 -11.580 15.765 -11.410 ;
        RECT 35.845 -11.580 36.015 -11.410 ;
        RECT 15.865 -18.960 16.035 -18.790 ;
        RECT 36.115 -18.960 36.285 -18.790 ;
      LAYER met1 ;
        RECT 13.440 6.710 35.115 7.135 ;
        RECT 14.840 4.935 15.970 5.255 ;
        RECT 35.260 4.935 36.220 5.255 ;
        RECT 13.440 -3.855 13.800 -3.685 ;
        RECT 15.915 -3.855 16.175 -2.035 ;
        RECT 13.440 -4.060 16.175 -3.855 ;
        RECT 33.690 -3.855 34.050 -3.685 ;
        RECT 36.165 -3.855 36.425 -2.035 ;
        RECT 33.690 -4.060 36.425 -3.855 ;
        RECT 14.820 -11.665 15.870 -11.345 ;
        RECT 34.935 -11.665 36.120 -11.345 ;
        RECT 13.340 -20.455 13.700 -20.285 ;
        RECT 15.815 -20.455 16.075 -18.635 ;
        RECT 13.340 -20.660 16.075 -20.455 ;
        RECT 33.590 -20.455 33.950 -20.285 ;
        RECT 36.065 -20.455 36.325 -18.635 ;
        RECT 33.590 -20.660 36.325 -20.455 ;
      LAYER via ;
        RECT 13.490 6.795 13.750 7.055 ;
        RECT 34.415 6.805 34.675 7.065 ;
        RECT 14.980 4.975 15.240 5.235 ;
        RECT 35.920 4.955 36.180 5.215 ;
        RECT 13.485 -3.995 13.745 -3.735 ;
        RECT 33.735 -3.995 33.995 -3.735 ;
        RECT 14.880 -11.625 15.140 -11.365 ;
        RECT 35.830 -11.645 36.090 -11.385 ;
        RECT 13.385 -20.595 13.645 -20.335 ;
        RECT 33.635 -20.595 33.895 -20.335 ;
      LAYER met2 ;
        RECT 13.435 8.075 15.250 9.855 ;
        RECT 13.440 -20.280 13.805 8.075 ;
        RECT 34.055 6.700 35.110 7.570 ;
        RECT 14.495 4.685 15.350 5.545 ;
        RECT 34.055 4.760 34.420 6.700 ;
        RECT 35.800 4.815 36.330 5.505 ;
        RECT 33.685 4.150 34.420 4.760 ;
        RECT 33.685 -3.680 34.055 4.150 ;
        RECT 14.395 -11.915 15.250 -11.055 ;
        RECT 33.690 -20.280 34.055 -3.680 ;
        RECT 35.460 -11.860 36.280 -11.235 ;
        RECT 13.340 -20.660 13.805 -20.280 ;
        RECT 33.590 -20.660 34.055 -20.280 ;
      LAYER via2 ;
        RECT 13.705 9.250 13.985 9.530 ;
        RECT 14.190 9.250 14.470 9.530 ;
        RECT 14.700 9.250 14.980 9.530 ;
        RECT 13.705 8.835 13.985 9.115 ;
        RECT 14.190 8.835 14.470 9.115 ;
        RECT 14.700 8.835 14.980 9.115 ;
        RECT 13.705 8.395 13.985 8.675 ;
        RECT 14.190 8.395 14.470 8.675 ;
        RECT 14.700 8.395 14.980 8.675 ;
        RECT 14.655 4.970 14.935 5.250 ;
        RECT 35.910 5.090 36.190 5.370 ;
        RECT 14.555 -11.630 14.835 -11.350 ;
        RECT 35.750 -11.735 36.030 -11.455 ;
      LAYER met3 ;
        RECT 13.435 8.075 15.250 9.855 ;
        RECT 14.495 5.465 15.350 5.545 ;
        RECT 14.495 4.975 36.275 5.465 ;
        RECT 14.495 4.685 15.350 4.975 ;
        RECT 14.395 -11.430 36.100 -11.055 ;
        RECT 14.395 -11.915 15.250 -11.430 ;
        RECT 35.680 -11.805 36.100 -11.430 ;
      LAYER via3 ;
        RECT 13.685 9.230 14.005 9.550 ;
        RECT 14.170 9.230 14.490 9.550 ;
        RECT 14.680 9.230 15.000 9.550 ;
        RECT 13.685 8.815 14.005 9.135 ;
        RECT 14.170 8.815 14.490 9.135 ;
        RECT 14.680 8.815 15.000 9.135 ;
        RECT 13.685 8.375 14.005 8.695 ;
        RECT 14.170 8.375 14.490 8.695 ;
        RECT 14.680 8.375 15.000 8.695 ;
        RECT 14.635 4.950 14.955 5.270 ;
        RECT 14.535 -11.650 14.855 -11.330 ;
      LAYER met4 ;
        RECT 13.510 -72.000 15.250 165.250 ;
    END
  END vccd1
  OBS
      LAYER pwell ;
        RECT 17.120 4.170 18.130 4.790 ;
        RECT 37.370 4.170 38.380 4.790 ;
        RECT -4.860 1.875 -3.850 2.495 ;
        RECT -3.645 1.235 -2.635 2.495 ;
        RECT -2.590 -0.765 -1.580 2.495 ;
        RECT -1.555 -4.775 -0.545 2.485 ;
        RECT 14.380 -4.595 15.390 2.665 ;
        RECT 17.015 0.340 17.635 0.910 ;
        RECT 16.985 -0.160 17.665 0.340 ;
        RECT 16.985 -0.670 17.895 -0.160 ;
        RECT 16.985 -1.180 17.665 -0.670 ;
        RECT 17.015 -1.750 17.635 -1.180 ;
        RECT 18.655 -4.595 19.665 2.665 ;
        RECT 34.630 -4.595 35.640 2.665 ;
        RECT 37.265 0.340 37.885 0.910 ;
        RECT 37.235 -0.160 37.915 0.340 ;
        RECT 37.235 -0.670 38.145 -0.160 ;
        RECT 37.235 -1.180 37.915 -0.670 ;
        RECT 37.265 -1.750 37.885 -1.180 ;
        RECT 38.905 -4.595 39.915 2.665 ;
        RECT 17.020 -12.430 18.030 -11.810 ;
        RECT 37.270 -12.430 38.280 -11.810 ;
        RECT 14.280 -21.195 15.290 -13.935 ;
        RECT 16.915 -16.260 17.535 -15.690 ;
        RECT 16.885 -16.760 17.565 -16.260 ;
        RECT 16.885 -17.270 17.795 -16.760 ;
        RECT 16.885 -17.780 17.565 -17.270 ;
        RECT 16.915 -18.350 17.535 -17.780 ;
        RECT 18.555 -21.195 19.565 -13.935 ;
        RECT 34.530 -21.195 35.540 -13.935 ;
        RECT 37.165 -16.260 37.785 -15.690 ;
        RECT 37.135 -16.760 37.815 -16.260 ;
        RECT 37.135 -17.270 38.045 -16.760 ;
        RECT 37.135 -17.780 37.815 -17.270 ;
        RECT 37.165 -18.350 37.785 -17.780 ;
        RECT 38.805 -21.195 39.815 -13.935 ;
      LAYER li1 ;
        RECT 16.195 4.940 16.365 5.270 ;
        RECT 36.445 4.940 36.615 5.270 ;
        RECT -4.190 2.020 -4.020 2.350 ;
        RECT -2.975 1.400 -2.805 2.350 ;
        RECT -1.920 -0.635 -1.750 2.350 ;
        RECT -0.885 -3.000 -0.715 2.350 ;
        RECT 15.050 -2.820 15.220 2.530 ;
        RECT 15.850 1.115 16.220 4.655 ;
        RECT 17.790 4.315 17.960 4.645 ;
        RECT 17.470 1.115 17.820 3.980 ;
        RECT 16.175 0.250 17.425 0.360 ;
        RECT 16.095 0.190 17.505 0.250 ;
        RECT 16.095 -0.080 16.495 0.190 ;
        RECT 15.895 -0.590 16.145 -0.260 ;
        RECT 16.325 -0.410 16.495 -0.080 ;
        RECT 16.675 -0.060 17.005 0.020 ;
        RECT 16.675 -0.230 17.085 -0.060 ;
        RECT 17.255 -0.080 17.505 0.190 ;
        RECT 16.915 -0.250 17.085 -0.230 ;
        RECT 16.325 -0.580 16.685 -0.410 ;
        RECT 16.915 -0.420 17.345 -0.250 ;
        RECT 16.515 -0.610 16.685 -0.580 ;
        RECT 16.095 -1.030 16.345 -0.760 ;
        RECT 16.515 -0.780 17.005 -0.610 ;
        RECT 16.675 -0.860 17.005 -0.780 ;
        RECT 17.175 -0.760 17.345 -0.420 ;
        RECT 17.515 -0.580 17.765 -0.250 ;
        RECT 17.175 -1.030 17.505 -0.760 ;
        RECT 16.095 -1.090 17.505 -1.030 ;
        RECT 16.175 -1.200 17.425 -1.090 ;
        RECT 19.325 -2.820 19.495 2.530 ;
        RECT 35.300 -2.820 35.470 2.530 ;
        RECT 36.100 1.115 36.470 4.655 ;
        RECT 38.040 4.315 38.210 4.645 ;
        RECT 37.720 1.115 38.070 3.980 ;
        RECT 36.425 0.250 37.675 0.360 ;
        RECT 36.345 0.190 37.755 0.250 ;
        RECT 36.345 -0.080 36.745 0.190 ;
        RECT 36.145 -0.590 36.395 -0.260 ;
        RECT 36.575 -0.410 36.745 -0.080 ;
        RECT 36.925 -0.060 37.255 0.020 ;
        RECT 36.925 -0.230 37.335 -0.060 ;
        RECT 37.505 -0.080 37.755 0.190 ;
        RECT 37.165 -0.250 37.335 -0.230 ;
        RECT 36.575 -0.580 36.935 -0.410 ;
        RECT 37.165 -0.420 37.595 -0.250 ;
        RECT 36.765 -0.610 36.935 -0.580 ;
        RECT 36.345 -1.030 36.595 -0.760 ;
        RECT 36.765 -0.780 37.255 -0.610 ;
        RECT 36.925 -0.860 37.255 -0.780 ;
        RECT 37.425 -0.760 37.595 -0.420 ;
        RECT 37.765 -0.580 38.015 -0.250 ;
        RECT 37.425 -1.030 37.755 -0.760 ;
        RECT 36.345 -1.090 37.755 -1.030 ;
        RECT 36.425 -1.200 37.675 -1.090 ;
        RECT 39.575 -2.820 39.745 2.530 ;
        RECT 16.095 -11.660 16.265 -11.330 ;
        RECT 36.345 -11.660 36.515 -11.330 ;
        RECT 14.950 -19.420 15.120 -14.070 ;
        RECT 15.750 -15.485 16.120 -11.945 ;
        RECT 17.690 -12.285 17.860 -11.955 ;
        RECT 17.370 -15.485 17.720 -12.620 ;
        RECT 16.075 -16.350 17.325 -16.240 ;
        RECT 15.995 -16.410 17.405 -16.350 ;
        RECT 15.995 -16.680 16.395 -16.410 ;
        RECT 15.795 -17.190 16.045 -16.860 ;
        RECT 16.225 -17.010 16.395 -16.680 ;
        RECT 16.575 -16.660 16.905 -16.580 ;
        RECT 16.575 -16.830 16.985 -16.660 ;
        RECT 17.155 -16.680 17.405 -16.410 ;
        RECT 16.815 -16.850 16.985 -16.830 ;
        RECT 16.225 -17.180 16.585 -17.010 ;
        RECT 16.815 -17.020 17.245 -16.850 ;
        RECT 16.415 -17.210 16.585 -17.180 ;
        RECT 15.995 -17.630 16.245 -17.360 ;
        RECT 16.415 -17.380 16.905 -17.210 ;
        RECT 16.575 -17.460 16.905 -17.380 ;
        RECT 17.075 -17.360 17.245 -17.020 ;
        RECT 17.415 -17.180 17.665 -16.850 ;
        RECT 17.075 -17.630 17.405 -17.360 ;
        RECT 15.995 -17.690 17.405 -17.630 ;
        RECT 16.075 -17.800 17.325 -17.690 ;
        RECT 19.225 -19.420 19.395 -14.070 ;
        RECT 35.200 -19.420 35.370 -14.070 ;
        RECT 36.000 -15.485 36.370 -11.945 ;
        RECT 37.940 -12.285 38.110 -11.955 ;
        RECT 37.620 -15.485 37.970 -12.620 ;
        RECT 36.325 -16.350 37.575 -16.240 ;
        RECT 36.245 -16.410 37.655 -16.350 ;
        RECT 36.245 -16.680 36.645 -16.410 ;
        RECT 36.045 -17.190 36.295 -16.860 ;
        RECT 36.475 -17.010 36.645 -16.680 ;
        RECT 36.825 -16.660 37.155 -16.580 ;
        RECT 36.825 -16.830 37.235 -16.660 ;
        RECT 37.405 -16.680 37.655 -16.410 ;
        RECT 37.065 -16.850 37.235 -16.830 ;
        RECT 36.475 -17.180 36.835 -17.010 ;
        RECT 37.065 -17.020 37.495 -16.850 ;
        RECT 36.665 -17.210 36.835 -17.180 ;
        RECT 36.245 -17.630 36.495 -17.360 ;
        RECT 36.665 -17.380 37.155 -17.210 ;
        RECT 36.825 -17.460 37.155 -17.380 ;
        RECT 37.325 -17.360 37.495 -17.020 ;
        RECT 37.665 -17.180 37.915 -16.850 ;
        RECT 37.325 -17.630 37.655 -17.360 ;
        RECT 36.245 -17.690 37.655 -17.630 ;
        RECT 36.325 -17.800 37.575 -17.690 ;
        RECT 39.475 -19.420 39.645 -14.070 ;
      LAYER mcon ;
        RECT 16.195 5.020 16.365 5.190 ;
        RECT 36.445 5.020 36.615 5.190 ;
        RECT 15.955 4.415 16.125 4.585 ;
        RECT -4.190 2.100 -4.020 2.270 ;
        RECT -2.975 1.975 -2.805 2.145 ;
        RECT -2.975 1.615 -2.805 1.785 ;
        RECT -1.920 1.800 -1.750 1.970 ;
        RECT -1.920 1.440 -1.750 1.610 ;
        RECT -1.920 1.080 -1.750 1.250 ;
        RECT -1.920 0.720 -1.750 0.890 ;
        RECT -1.920 0.360 -1.750 0.530 ;
        RECT -1.920 0.000 -1.750 0.170 ;
        RECT -1.920 -0.360 -1.750 -0.190 ;
        RECT -0.885 1.960 -0.715 2.130 ;
        RECT -0.885 1.600 -0.715 1.770 ;
        RECT -0.885 1.240 -0.715 1.410 ;
        RECT -0.885 0.880 -0.715 1.050 ;
        RECT -0.885 0.520 -0.715 0.690 ;
        RECT -0.885 0.160 -0.715 0.330 ;
        RECT -0.885 -0.200 -0.715 -0.030 ;
        RECT -0.885 -0.560 -0.715 -0.390 ;
        RECT -0.885 -0.920 -0.715 -0.750 ;
        RECT -0.885 -1.280 -0.715 -1.110 ;
        RECT -0.885 -1.640 -0.715 -1.470 ;
        RECT -0.885 -2.000 -0.715 -1.830 ;
        RECT -0.885 -2.360 -0.715 -2.190 ;
        RECT -0.885 -2.720 -0.715 -2.550 ;
        RECT 15.050 2.140 15.220 2.310 ;
        RECT 15.050 1.780 15.220 1.950 ;
        RECT 15.050 1.420 15.220 1.590 ;
        RECT 15.050 1.060 15.220 1.230 ;
        RECT 17.790 4.395 17.960 4.565 ;
        RECT 36.205 4.395 36.375 4.565 ;
        RECT 15.950 1.225 16.120 1.395 ;
        RECT 17.550 3.760 17.720 3.930 ;
        RECT 17.535 1.220 17.705 1.390 ;
        RECT 19.325 2.140 19.495 2.310 ;
        RECT 19.325 1.780 19.495 1.950 ;
        RECT 19.325 1.420 19.495 1.590 ;
        RECT 15.050 0.700 15.220 0.870 ;
        RECT 15.050 0.340 15.220 0.510 ;
        RECT 19.325 1.060 19.495 1.230 ;
        RECT 19.325 0.700 19.495 0.870 ;
        RECT 19.325 0.340 19.495 0.510 ;
        RECT 15.050 -0.020 15.220 0.150 ;
        RECT 15.050 -0.380 15.220 -0.210 ;
        RECT 15.050 -0.740 15.220 -0.570 ;
        RECT 15.975 -0.510 16.145 -0.340 ;
        RECT 19.325 -0.020 19.495 0.150 ;
        RECT 15.050 -1.100 15.220 -0.930 ;
        RECT 17.515 -0.500 17.685 -0.330 ;
        RECT 19.325 -0.380 19.495 -0.210 ;
        RECT 19.325 -0.740 19.495 -0.570 ;
        RECT 19.325 -1.100 19.495 -0.930 ;
        RECT 15.050 -1.460 15.220 -1.290 ;
        RECT 15.050 -1.820 15.220 -1.650 ;
        RECT 15.050 -2.180 15.220 -2.010 ;
        RECT 15.050 -2.540 15.220 -2.370 ;
        RECT 19.325 -1.460 19.495 -1.290 ;
        RECT 19.325 -1.820 19.495 -1.650 ;
        RECT 19.325 -2.180 19.495 -2.010 ;
        RECT 19.325 -2.540 19.495 -2.370 ;
        RECT 35.300 2.140 35.470 2.310 ;
        RECT 35.300 1.780 35.470 1.950 ;
        RECT 35.300 1.420 35.470 1.590 ;
        RECT 35.300 1.060 35.470 1.230 ;
        RECT 38.040 4.395 38.210 4.565 ;
        RECT 36.200 1.225 36.370 1.395 ;
        RECT 37.800 3.755 37.970 3.925 ;
        RECT 37.785 1.220 37.955 1.390 ;
        RECT 39.575 2.140 39.745 2.310 ;
        RECT 39.575 1.780 39.745 1.950 ;
        RECT 39.575 1.420 39.745 1.590 ;
        RECT 35.300 0.700 35.470 0.870 ;
        RECT 35.300 0.340 35.470 0.510 ;
        RECT 39.575 1.060 39.745 1.230 ;
        RECT 39.575 0.700 39.745 0.870 ;
        RECT 39.575 0.340 39.745 0.510 ;
        RECT 35.300 -0.020 35.470 0.150 ;
        RECT 35.300 -0.380 35.470 -0.210 ;
        RECT 35.300 -0.740 35.470 -0.570 ;
        RECT 36.225 -0.510 36.395 -0.340 ;
        RECT 39.575 -0.020 39.745 0.150 ;
        RECT 35.300 -1.100 35.470 -0.930 ;
        RECT 37.765 -0.500 37.935 -0.330 ;
        RECT 39.575 -0.380 39.745 -0.210 ;
        RECT 39.575 -0.740 39.745 -0.570 ;
        RECT 39.575 -1.100 39.745 -0.930 ;
        RECT 35.300 -1.460 35.470 -1.290 ;
        RECT 35.300 -1.820 35.470 -1.650 ;
        RECT 35.300 -2.180 35.470 -2.010 ;
        RECT 35.300 -2.540 35.470 -2.370 ;
        RECT 39.575 -1.460 39.745 -1.290 ;
        RECT 39.575 -1.820 39.745 -1.650 ;
        RECT 39.575 -2.180 39.745 -2.010 ;
        RECT 39.575 -2.540 39.745 -2.370 ;
        RECT 16.095 -11.580 16.265 -11.410 ;
        RECT 36.345 -11.580 36.515 -11.410 ;
        RECT 15.855 -12.185 16.025 -12.015 ;
        RECT 14.950 -14.460 15.120 -14.290 ;
        RECT 14.950 -14.820 15.120 -14.650 ;
        RECT 14.950 -15.180 15.120 -15.010 ;
        RECT 14.950 -15.540 15.120 -15.370 ;
        RECT 17.690 -12.205 17.860 -12.035 ;
        RECT 36.105 -12.190 36.275 -12.020 ;
        RECT 15.850 -15.375 16.020 -15.205 ;
        RECT 17.450 -12.840 17.620 -12.670 ;
        RECT 17.435 -15.380 17.605 -15.210 ;
        RECT 19.225 -14.460 19.395 -14.290 ;
        RECT 19.225 -14.820 19.395 -14.650 ;
        RECT 19.225 -15.180 19.395 -15.010 ;
        RECT 14.950 -15.900 15.120 -15.730 ;
        RECT 14.950 -16.260 15.120 -16.090 ;
        RECT 19.225 -15.540 19.395 -15.370 ;
        RECT 19.225 -15.900 19.395 -15.730 ;
        RECT 19.225 -16.260 19.395 -16.090 ;
        RECT 14.950 -16.620 15.120 -16.450 ;
        RECT 14.950 -16.980 15.120 -16.810 ;
        RECT 14.950 -17.340 15.120 -17.170 ;
        RECT 15.875 -17.110 16.045 -16.940 ;
        RECT 19.225 -16.620 19.395 -16.450 ;
        RECT 14.950 -17.700 15.120 -17.530 ;
        RECT 17.415 -17.100 17.585 -16.930 ;
        RECT 19.225 -16.980 19.395 -16.810 ;
        RECT 19.225 -17.340 19.395 -17.170 ;
        RECT 19.225 -17.700 19.395 -17.530 ;
        RECT 14.950 -18.060 15.120 -17.890 ;
        RECT 14.950 -18.420 15.120 -18.250 ;
        RECT 14.950 -18.780 15.120 -18.610 ;
        RECT 14.950 -19.140 15.120 -18.970 ;
        RECT 19.225 -18.060 19.395 -17.890 ;
        RECT 19.225 -18.420 19.395 -18.250 ;
        RECT 19.225 -18.780 19.395 -18.610 ;
        RECT 19.225 -19.140 19.395 -18.970 ;
        RECT 35.200 -14.460 35.370 -14.290 ;
        RECT 35.200 -14.820 35.370 -14.650 ;
        RECT 35.200 -15.180 35.370 -15.010 ;
        RECT 35.200 -15.540 35.370 -15.370 ;
        RECT 37.940 -12.205 38.110 -12.035 ;
        RECT 36.100 -15.375 36.270 -15.205 ;
        RECT 37.700 -12.840 37.870 -12.670 ;
        RECT 37.685 -15.380 37.855 -15.210 ;
        RECT 39.475 -14.460 39.645 -14.290 ;
        RECT 39.475 -14.820 39.645 -14.650 ;
        RECT 39.475 -15.180 39.645 -15.010 ;
        RECT 35.200 -15.900 35.370 -15.730 ;
        RECT 35.200 -16.260 35.370 -16.090 ;
        RECT 39.475 -15.540 39.645 -15.370 ;
        RECT 39.475 -15.900 39.645 -15.730 ;
        RECT 39.475 -16.260 39.645 -16.090 ;
        RECT 35.200 -16.620 35.370 -16.450 ;
        RECT 35.200 -16.980 35.370 -16.810 ;
        RECT 35.200 -17.340 35.370 -17.170 ;
        RECT 36.125 -17.110 36.295 -16.940 ;
        RECT 39.475 -16.620 39.645 -16.450 ;
        RECT 35.200 -17.700 35.370 -17.530 ;
        RECT 37.665 -17.100 37.835 -16.930 ;
        RECT 39.475 -16.980 39.645 -16.810 ;
        RECT 39.475 -17.340 39.645 -17.170 ;
        RECT 39.475 -17.700 39.645 -17.530 ;
        RECT 35.200 -18.060 35.370 -17.890 ;
        RECT 35.200 -18.420 35.370 -18.250 ;
        RECT 35.200 -18.780 35.370 -18.610 ;
        RECT 35.200 -19.140 35.370 -18.970 ;
        RECT 39.475 -18.060 39.645 -17.890 ;
        RECT 39.475 -18.420 39.645 -18.250 ;
        RECT 39.475 -18.780 39.645 -18.610 ;
        RECT 39.475 -19.140 39.645 -18.970 ;
      LAYER met1 ;
        RECT 16.165 4.960 16.395 5.270 ;
        RECT 36.415 4.960 36.645 5.270 ;
        RECT 16.210 4.795 16.350 4.960 ;
        RECT 36.460 4.795 36.600 4.960 ;
        RECT 15.955 4.655 16.350 4.795 ;
        RECT 36.205 4.655 36.600 4.795 ;
        RECT 15.850 4.265 16.220 4.655 ;
        RECT 17.760 4.335 17.990 4.645 ;
        RECT 17.805 4.170 17.945 4.335 ;
        RECT 36.100 4.275 36.470 4.655 ;
        RECT 38.010 4.335 38.240 4.645 ;
        RECT 38.055 4.170 38.195 4.335 ;
        RECT 17.550 4.030 17.945 4.170 ;
        RECT 37.800 4.030 38.195 4.170 ;
        RECT 17.470 3.670 17.820 4.030 ;
        RECT 37.720 3.670 38.070 4.030 ;
        RECT -4.530 2.950 -4.210 3.210 ;
        RECT -3.315 2.950 -2.995 3.210 ;
        RECT -2.260 2.950 -1.940 3.210 ;
        RECT -1.225 2.950 -0.905 3.210 ;
        RECT 14.710 3.130 15.030 3.390 ;
        RECT 18.985 3.130 19.305 3.390 ;
        RECT 34.960 3.130 35.280 3.390 ;
        RECT 39.235 3.130 39.555 3.390 ;
        RECT -4.430 2.635 -4.270 2.950 ;
        RECT -3.215 2.635 -3.055 2.950 ;
        RECT -2.160 2.635 -2.000 2.950 ;
        RECT -1.125 2.635 -0.965 2.950 ;
        RECT 14.810 2.815 14.970 3.130 ;
        RECT 19.085 2.815 19.245 3.130 ;
        RECT 35.060 2.815 35.220 3.130 ;
        RECT 39.335 2.815 39.495 3.130 ;
        RECT 14.810 2.675 15.205 2.815 ;
        RECT 19.085 2.675 19.480 2.815 ;
        RECT 35.060 2.675 35.455 2.815 ;
        RECT 39.335 2.675 39.730 2.815 ;
        RECT -4.430 2.495 -4.035 2.635 ;
        RECT -3.215 2.495 -2.820 2.635 ;
        RECT -2.160 2.495 -1.765 2.635 ;
        RECT -1.125 2.495 -0.730 2.635 ;
        RECT 15.065 2.510 15.205 2.675 ;
        RECT 19.340 2.510 19.480 2.675 ;
        RECT 35.315 2.510 35.455 2.675 ;
        RECT 39.590 2.510 39.730 2.675 ;
        RECT -4.175 2.330 -4.035 2.495 ;
        RECT -2.960 2.330 -2.820 2.495 ;
        RECT -1.905 2.330 -1.765 2.495 ;
        RECT -0.870 2.330 -0.730 2.495 ;
        RECT -4.220 2.020 -3.990 2.330 ;
        RECT -3.005 1.395 -2.775 2.330 ;
        RECT -1.950 -0.635 -1.720 2.330 ;
        RECT -0.915 -3.000 -0.685 2.330 ;
        RECT 15.020 -2.820 15.250 2.510 ;
        RECT 15.915 0.360 16.175 1.490 ;
        RECT 17.505 0.780 17.745 1.490 ;
        RECT 15.915 0.040 16.235 0.360 ;
        RECT 15.915 -0.280 16.175 0.040 ;
        RECT 17.485 -0.260 17.745 0.780 ;
        RECT 15.915 -0.570 16.205 -0.280 ;
        RECT 15.915 -1.620 16.175 -0.570 ;
        RECT 17.425 -0.580 17.745 -0.260 ;
        RECT 17.485 -1.620 17.745 -0.580 ;
        RECT 19.295 -2.820 19.525 2.510 ;
        RECT 35.270 -2.820 35.500 2.510 ;
        RECT 36.165 0.360 36.425 1.490 ;
        RECT 37.755 0.780 37.995 1.490 ;
        RECT 36.165 0.040 36.485 0.360 ;
        RECT 36.165 -0.280 36.425 0.040 ;
        RECT 37.735 -0.260 37.995 0.780 ;
        RECT 36.165 -0.570 36.455 -0.280 ;
        RECT 36.165 -1.620 36.425 -0.570 ;
        RECT 37.675 -0.580 37.995 -0.260 ;
        RECT 37.735 -1.620 37.995 -0.580 ;
        RECT 39.545 -2.820 39.775 2.510 ;
        RECT 16.065 -11.640 16.295 -11.330 ;
        RECT 36.315 -11.640 36.545 -11.330 ;
        RECT 16.110 -11.805 16.250 -11.640 ;
        RECT 36.360 -11.805 36.500 -11.640 ;
        RECT 15.855 -11.945 16.250 -11.805 ;
        RECT 36.105 -11.945 36.500 -11.805 ;
        RECT 15.750 -12.295 16.120 -11.945 ;
        RECT 17.660 -12.265 17.890 -11.955 ;
        RECT 17.705 -12.430 17.845 -12.265 ;
        RECT 36.000 -12.275 36.370 -11.945 ;
        RECT 37.910 -12.265 38.140 -11.955 ;
        RECT 37.955 -12.430 38.095 -12.265 ;
        RECT 17.450 -12.570 17.845 -12.430 ;
        RECT 37.700 -12.570 38.095 -12.430 ;
        RECT 17.370 -12.985 17.720 -12.570 ;
        RECT 37.620 -12.920 37.970 -12.570 ;
        RECT 14.610 -13.470 14.930 -13.210 ;
        RECT 18.885 -13.470 19.205 -13.210 ;
        RECT 34.860 -13.470 35.180 -13.210 ;
        RECT 39.135 -13.470 39.455 -13.210 ;
        RECT 14.710 -13.785 14.870 -13.470 ;
        RECT 18.985 -13.785 19.145 -13.470 ;
        RECT 34.960 -13.785 35.120 -13.470 ;
        RECT 39.235 -13.785 39.395 -13.470 ;
        RECT 14.710 -13.925 15.105 -13.785 ;
        RECT 18.985 -13.925 19.380 -13.785 ;
        RECT 34.960 -13.925 35.355 -13.785 ;
        RECT 39.235 -13.925 39.630 -13.785 ;
        RECT 14.965 -14.090 15.105 -13.925 ;
        RECT 19.240 -14.090 19.380 -13.925 ;
        RECT 35.215 -14.090 35.355 -13.925 ;
        RECT 39.490 -14.090 39.630 -13.925 ;
        RECT 14.920 -19.420 15.150 -14.090 ;
        RECT 15.815 -16.240 16.075 -15.110 ;
        RECT 17.405 -15.820 17.645 -15.110 ;
        RECT 15.815 -16.560 16.135 -16.240 ;
        RECT 15.815 -16.880 16.075 -16.560 ;
        RECT 17.385 -16.860 17.645 -15.820 ;
        RECT 15.815 -17.170 16.105 -16.880 ;
        RECT 15.815 -18.220 16.075 -17.170 ;
        RECT 17.325 -17.180 17.645 -16.860 ;
        RECT 17.385 -18.220 17.645 -17.180 ;
        RECT 19.195 -19.420 19.425 -14.090 ;
        RECT 35.170 -19.420 35.400 -14.090 ;
        RECT 36.065 -16.240 36.325 -15.110 ;
        RECT 37.655 -15.820 37.895 -15.110 ;
        RECT 36.065 -16.560 36.385 -16.240 ;
        RECT 36.065 -16.880 36.325 -16.560 ;
        RECT 37.635 -16.860 37.895 -15.820 ;
        RECT 36.065 -17.170 36.355 -16.880 ;
        RECT 36.065 -18.220 36.325 -17.170 ;
        RECT 37.575 -17.180 37.895 -16.860 ;
        RECT 37.635 -18.220 37.895 -17.180 ;
        RECT 39.445 -19.420 39.675 -14.090 ;
      LAYER via ;
        RECT 15.945 0.070 16.205 0.330 ;
        RECT 17.455 -0.550 17.715 -0.290 ;
        RECT 36.195 0.070 36.455 0.330 ;
        RECT 37.705 -0.550 37.965 -0.290 ;
        RECT 15.845 -16.530 16.105 -16.270 ;
        RECT 17.355 -17.150 17.615 -16.890 ;
        RECT 36.095 -16.530 36.355 -16.270 ;
        RECT 37.605 -17.150 37.865 -16.890 ;
      LAYER met2 ;
        RECT 15.895 0.040 17.765 0.360 ;
        RECT 36.145 0.040 38.015 0.360 ;
        RECT 15.895 -0.580 17.765 -0.260 ;
        RECT 36.145 -0.580 38.015 -0.260 ;
        RECT 15.895 -1.200 17.765 -0.880 ;
        RECT 36.145 -1.200 38.015 -0.880 ;
        RECT 15.795 -16.560 17.665 -16.240 ;
        RECT 36.045 -16.560 37.915 -16.240 ;
        RECT 15.795 -17.180 17.665 -16.860 ;
        RECT 36.045 -17.180 37.915 -16.860 ;
        RECT 15.795 -17.800 17.665 -17.480 ;
        RECT 36.045 -17.800 37.915 -17.480 ;
  END
END rram_test
END LIBRARY


magic
tech sky130B
magscale 1 2
timestamp 1671441199
<< obsli1 >>
rect 1104 2159 582820 701777
<< obsm1 >>
rect 566 1708 583450 701808
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< obsm2 >>
rect 572 703464 8030 703610
rect 8254 703464 24222 703610
rect 24446 703464 40414 703610
rect 40638 703464 56698 703610
rect 56922 703464 72890 703610
rect 73114 703464 89082 703610
rect 89306 703464 105366 703610
rect 105590 703464 121558 703610
rect 121782 703464 137750 703610
rect 137974 703464 154034 703610
rect 154258 703464 170226 703610
rect 170450 703464 186418 703610
rect 186642 703464 202702 703610
rect 202926 703464 218894 703610
rect 219118 703464 235086 703610
rect 235310 703464 251370 703610
rect 251594 703464 267562 703610
rect 267786 703464 283754 703610
rect 283978 703464 300038 703610
rect 300262 703464 316230 703610
rect 316454 703464 332422 703610
rect 332646 703464 348706 703610
rect 348930 703464 364898 703610
rect 365122 703464 381090 703610
rect 381314 703464 397374 703610
rect 397598 703464 413566 703610
rect 413790 703464 429758 703610
rect 429982 703464 446042 703610
rect 446266 703464 462234 703610
rect 462458 703464 478426 703610
rect 478650 703464 494710 703610
rect 494934 703464 510902 703610
rect 511126 703464 527094 703610
rect 527318 703464 543378 703610
rect 543602 703464 559570 703610
rect 559794 703464 575762 703610
rect 575986 703464 583444 703610
rect 572 536 583444 703464
rect 710 190 1590 536
rect 1814 190 2786 536
rect 3010 190 3982 536
rect 4206 190 5178 536
rect 5402 190 6374 536
rect 6598 190 7570 536
rect 7794 190 8674 536
rect 8898 190 9870 536
rect 10094 190 11066 536
rect 11290 190 12262 536
rect 12486 190 13458 536
rect 13682 190 14654 536
rect 14878 190 15850 536
rect 16074 190 16954 536
rect 17178 190 18150 536
rect 18374 190 19346 536
rect 19570 190 20542 536
rect 20766 190 21738 536
rect 21962 190 22934 536
rect 23158 190 24130 536
rect 24354 190 25234 536
rect 25458 190 26430 536
rect 26654 190 27626 536
rect 27850 190 28822 536
rect 29046 190 30018 536
rect 30242 190 31214 536
rect 31438 190 32318 536
rect 32542 190 33514 536
rect 33738 190 34710 536
rect 34934 190 35906 536
rect 36130 190 37102 536
rect 37326 190 38298 536
rect 38522 190 39494 536
rect 39718 190 40598 536
rect 40822 190 41794 536
rect 42018 190 42990 536
rect 43214 190 44186 536
rect 44410 190 45382 536
rect 45606 190 46578 536
rect 46802 190 47774 536
rect 47998 190 48878 536
rect 49102 190 50074 536
rect 50298 190 51270 536
rect 51494 190 52466 536
rect 52690 190 53662 536
rect 53886 190 54858 536
rect 55082 190 55962 536
rect 56186 190 57158 536
rect 57382 190 58354 536
rect 58578 190 59550 536
rect 59774 190 60746 536
rect 60970 190 61942 536
rect 62166 190 63138 536
rect 63362 190 64242 536
rect 64466 190 65438 536
rect 65662 190 66634 536
rect 66858 190 67830 536
rect 68054 190 69026 536
rect 69250 190 70222 536
rect 70446 190 71418 536
rect 71642 190 72522 536
rect 72746 190 73718 536
rect 73942 190 74914 536
rect 75138 190 76110 536
rect 76334 190 77306 536
rect 77530 190 78502 536
rect 78726 190 79606 536
rect 79830 190 80802 536
rect 81026 190 81998 536
rect 82222 190 83194 536
rect 83418 190 84390 536
rect 84614 190 85586 536
rect 85810 190 86782 536
rect 87006 190 87886 536
rect 88110 190 89082 536
rect 89306 190 90278 536
rect 90502 190 91474 536
rect 91698 190 92670 536
rect 92894 190 93866 536
rect 94090 190 95062 536
rect 95286 190 96166 536
rect 96390 190 97362 536
rect 97586 190 98558 536
rect 98782 190 99754 536
rect 99978 190 100950 536
rect 101174 190 102146 536
rect 102370 190 103250 536
rect 103474 190 104446 536
rect 104670 190 105642 536
rect 105866 190 106838 536
rect 107062 190 108034 536
rect 108258 190 109230 536
rect 109454 190 110426 536
rect 110650 190 111530 536
rect 111754 190 112726 536
rect 112950 190 113922 536
rect 114146 190 115118 536
rect 115342 190 116314 536
rect 116538 190 117510 536
rect 117734 190 118706 536
rect 118930 190 119810 536
rect 120034 190 121006 536
rect 121230 190 122202 536
rect 122426 190 123398 536
rect 123622 190 124594 536
rect 124818 190 125790 536
rect 126014 190 126894 536
rect 127118 190 128090 536
rect 128314 190 129286 536
rect 129510 190 130482 536
rect 130706 190 131678 536
rect 131902 190 132874 536
rect 133098 190 134070 536
rect 134294 190 135174 536
rect 135398 190 136370 536
rect 136594 190 137566 536
rect 137790 190 138762 536
rect 138986 190 139958 536
rect 140182 190 141154 536
rect 141378 190 142350 536
rect 142574 190 143454 536
rect 143678 190 144650 536
rect 144874 190 145846 536
rect 146070 190 147042 536
rect 147266 190 148238 536
rect 148462 190 149434 536
rect 149658 190 150538 536
rect 150762 190 151734 536
rect 151958 190 152930 536
rect 153154 190 154126 536
rect 154350 190 155322 536
rect 155546 190 156518 536
rect 156742 190 157714 536
rect 157938 190 158818 536
rect 159042 190 160014 536
rect 160238 190 161210 536
rect 161434 190 162406 536
rect 162630 190 163602 536
rect 163826 190 164798 536
rect 165022 190 165994 536
rect 166218 190 167098 536
rect 167322 190 168294 536
rect 168518 190 169490 536
rect 169714 190 170686 536
rect 170910 190 171882 536
rect 172106 190 173078 536
rect 173302 190 174182 536
rect 174406 190 175378 536
rect 175602 190 176574 536
rect 176798 190 177770 536
rect 177994 190 178966 536
rect 179190 190 180162 536
rect 180386 190 181358 536
rect 181582 190 182462 536
rect 182686 190 183658 536
rect 183882 190 184854 536
rect 185078 190 186050 536
rect 186274 190 187246 536
rect 187470 190 188442 536
rect 188666 190 189638 536
rect 189862 190 190742 536
rect 190966 190 191938 536
rect 192162 190 193134 536
rect 193358 190 194330 536
rect 194554 190 195526 536
rect 195750 190 196722 536
rect 196946 190 197826 536
rect 198050 190 199022 536
rect 199246 190 200218 536
rect 200442 190 201414 536
rect 201638 190 202610 536
rect 202834 190 203806 536
rect 204030 190 205002 536
rect 205226 190 206106 536
rect 206330 190 207302 536
rect 207526 190 208498 536
rect 208722 190 209694 536
rect 209918 190 210890 536
rect 211114 190 212086 536
rect 212310 190 213282 536
rect 213506 190 214386 536
rect 214610 190 215582 536
rect 215806 190 216778 536
rect 217002 190 217974 536
rect 218198 190 219170 536
rect 219394 190 220366 536
rect 220590 190 221470 536
rect 221694 190 222666 536
rect 222890 190 223862 536
rect 224086 190 225058 536
rect 225282 190 226254 536
rect 226478 190 227450 536
rect 227674 190 228646 536
rect 228870 190 229750 536
rect 229974 190 230946 536
rect 231170 190 232142 536
rect 232366 190 233338 536
rect 233562 190 234534 536
rect 234758 190 235730 536
rect 235954 190 236926 536
rect 237150 190 238030 536
rect 238254 190 239226 536
rect 239450 190 240422 536
rect 240646 190 241618 536
rect 241842 190 242814 536
rect 243038 190 244010 536
rect 244234 190 245114 536
rect 245338 190 246310 536
rect 246534 190 247506 536
rect 247730 190 248702 536
rect 248926 190 249898 536
rect 250122 190 251094 536
rect 251318 190 252290 536
rect 252514 190 253394 536
rect 253618 190 254590 536
rect 254814 190 255786 536
rect 256010 190 256982 536
rect 257206 190 258178 536
rect 258402 190 259374 536
rect 259598 190 260570 536
rect 260794 190 261674 536
rect 261898 190 262870 536
rect 263094 190 264066 536
rect 264290 190 265262 536
rect 265486 190 266458 536
rect 266682 190 267654 536
rect 267878 190 268758 536
rect 268982 190 269954 536
rect 270178 190 271150 536
rect 271374 190 272346 536
rect 272570 190 273542 536
rect 273766 190 274738 536
rect 274962 190 275934 536
rect 276158 190 277038 536
rect 277262 190 278234 536
rect 278458 190 279430 536
rect 279654 190 280626 536
rect 280850 190 281822 536
rect 282046 190 283018 536
rect 283242 190 284214 536
rect 284438 190 285318 536
rect 285542 190 286514 536
rect 286738 190 287710 536
rect 287934 190 288906 536
rect 289130 190 290102 536
rect 290326 190 291298 536
rect 291522 190 292494 536
rect 292718 190 293598 536
rect 293822 190 294794 536
rect 295018 190 295990 536
rect 296214 190 297186 536
rect 297410 190 298382 536
rect 298606 190 299578 536
rect 299802 190 300682 536
rect 300906 190 301878 536
rect 302102 190 303074 536
rect 303298 190 304270 536
rect 304494 190 305466 536
rect 305690 190 306662 536
rect 306886 190 307858 536
rect 308082 190 308962 536
rect 309186 190 310158 536
rect 310382 190 311354 536
rect 311578 190 312550 536
rect 312774 190 313746 536
rect 313970 190 314942 536
rect 315166 190 316138 536
rect 316362 190 317242 536
rect 317466 190 318438 536
rect 318662 190 319634 536
rect 319858 190 320830 536
rect 321054 190 322026 536
rect 322250 190 323222 536
rect 323446 190 324326 536
rect 324550 190 325522 536
rect 325746 190 326718 536
rect 326942 190 327914 536
rect 328138 190 329110 536
rect 329334 190 330306 536
rect 330530 190 331502 536
rect 331726 190 332606 536
rect 332830 190 333802 536
rect 334026 190 334998 536
rect 335222 190 336194 536
rect 336418 190 337390 536
rect 337614 190 338586 536
rect 338810 190 339782 536
rect 340006 190 340886 536
rect 341110 190 342082 536
rect 342306 190 343278 536
rect 343502 190 344474 536
rect 344698 190 345670 536
rect 345894 190 346866 536
rect 347090 190 347970 536
rect 348194 190 349166 536
rect 349390 190 350362 536
rect 350586 190 351558 536
rect 351782 190 352754 536
rect 352978 190 353950 536
rect 354174 190 355146 536
rect 355370 190 356250 536
rect 356474 190 357446 536
rect 357670 190 358642 536
rect 358866 190 359838 536
rect 360062 190 361034 536
rect 361258 190 362230 536
rect 362454 190 363426 536
rect 363650 190 364530 536
rect 364754 190 365726 536
rect 365950 190 366922 536
rect 367146 190 368118 536
rect 368342 190 369314 536
rect 369538 190 370510 536
rect 370734 190 371614 536
rect 371838 190 372810 536
rect 373034 190 374006 536
rect 374230 190 375202 536
rect 375426 190 376398 536
rect 376622 190 377594 536
rect 377818 190 378790 536
rect 379014 190 379894 536
rect 380118 190 381090 536
rect 381314 190 382286 536
rect 382510 190 383482 536
rect 383706 190 384678 536
rect 384902 190 385874 536
rect 386098 190 387070 536
rect 387294 190 388174 536
rect 388398 190 389370 536
rect 389594 190 390566 536
rect 390790 190 391762 536
rect 391986 190 392958 536
rect 393182 190 394154 536
rect 394378 190 395258 536
rect 395482 190 396454 536
rect 396678 190 397650 536
rect 397874 190 398846 536
rect 399070 190 400042 536
rect 400266 190 401238 536
rect 401462 190 402434 536
rect 402658 190 403538 536
rect 403762 190 404734 536
rect 404958 190 405930 536
rect 406154 190 407126 536
rect 407350 190 408322 536
rect 408546 190 409518 536
rect 409742 190 410714 536
rect 410938 190 411818 536
rect 412042 190 413014 536
rect 413238 190 414210 536
rect 414434 190 415406 536
rect 415630 190 416602 536
rect 416826 190 417798 536
rect 418022 190 418902 536
rect 419126 190 420098 536
rect 420322 190 421294 536
rect 421518 190 422490 536
rect 422714 190 423686 536
rect 423910 190 424882 536
rect 425106 190 426078 536
rect 426302 190 427182 536
rect 427406 190 428378 536
rect 428602 190 429574 536
rect 429798 190 430770 536
rect 430994 190 431966 536
rect 432190 190 433162 536
rect 433386 190 434358 536
rect 434582 190 435462 536
rect 435686 190 436658 536
rect 436882 190 437854 536
rect 438078 190 439050 536
rect 439274 190 440246 536
rect 440470 190 441442 536
rect 441666 190 442546 536
rect 442770 190 443742 536
rect 443966 190 444938 536
rect 445162 190 446134 536
rect 446358 190 447330 536
rect 447554 190 448526 536
rect 448750 190 449722 536
rect 449946 190 450826 536
rect 451050 190 452022 536
rect 452246 190 453218 536
rect 453442 190 454414 536
rect 454638 190 455610 536
rect 455834 190 456806 536
rect 457030 190 458002 536
rect 458226 190 459106 536
rect 459330 190 460302 536
rect 460526 190 461498 536
rect 461722 190 462694 536
rect 462918 190 463890 536
rect 464114 190 465086 536
rect 465310 190 466190 536
rect 466414 190 467386 536
rect 467610 190 468582 536
rect 468806 190 469778 536
rect 470002 190 470974 536
rect 471198 190 472170 536
rect 472394 190 473366 536
rect 473590 190 474470 536
rect 474694 190 475666 536
rect 475890 190 476862 536
rect 477086 190 478058 536
rect 478282 190 479254 536
rect 479478 190 480450 536
rect 480674 190 481646 536
rect 481870 190 482750 536
rect 482974 190 483946 536
rect 484170 190 485142 536
rect 485366 190 486338 536
rect 486562 190 487534 536
rect 487758 190 488730 536
rect 488954 190 489834 536
rect 490058 190 491030 536
rect 491254 190 492226 536
rect 492450 190 493422 536
rect 493646 190 494618 536
rect 494842 190 495814 536
rect 496038 190 497010 536
rect 497234 190 498114 536
rect 498338 190 499310 536
rect 499534 190 500506 536
rect 500730 190 501702 536
rect 501926 190 502898 536
rect 503122 190 504094 536
rect 504318 190 505290 536
rect 505514 190 506394 536
rect 506618 190 507590 536
rect 507814 190 508786 536
rect 509010 190 509982 536
rect 510206 190 511178 536
rect 511402 190 512374 536
rect 512598 190 513478 536
rect 513702 190 514674 536
rect 514898 190 515870 536
rect 516094 190 517066 536
rect 517290 190 518262 536
rect 518486 190 519458 536
rect 519682 190 520654 536
rect 520878 190 521758 536
rect 521982 190 522954 536
rect 523178 190 524150 536
rect 524374 190 525346 536
rect 525570 190 526542 536
rect 526766 190 527738 536
rect 527962 190 528934 536
rect 529158 190 530038 536
rect 530262 190 531234 536
rect 531458 190 532430 536
rect 532654 190 533626 536
rect 533850 190 534822 536
rect 535046 190 536018 536
rect 536242 190 537122 536
rect 537346 190 538318 536
rect 538542 190 539514 536
rect 539738 190 540710 536
rect 540934 190 541906 536
rect 542130 190 543102 536
rect 543326 190 544298 536
rect 544522 190 545402 536
rect 545626 190 546598 536
rect 546822 190 547794 536
rect 548018 190 548990 536
rect 549214 190 550186 536
rect 550410 190 551382 536
rect 551606 190 552578 536
rect 552802 190 553682 536
rect 553906 190 554878 536
rect 555102 190 556074 536
rect 556298 190 557270 536
rect 557494 190 558466 536
rect 558690 190 559662 536
rect 559886 190 560766 536
rect 560990 190 561962 536
rect 562186 190 563158 536
rect 563382 190 564354 536
rect 564578 190 565550 536
rect 565774 190 566746 536
rect 566970 190 567942 536
rect 568166 190 569046 536
rect 569270 190 570242 536
rect 570466 190 571438 536
rect 571662 190 572634 536
rect 572858 190 573830 536
rect 574054 190 575026 536
rect 575250 190 576222 536
rect 576446 190 577326 536
rect 577550 190 578522 536
rect 578746 190 579718 536
rect 579942 190 580914 536
rect 581138 190 582110 536
rect 582334 190 583306 536
<< metal3 >>
rect -960 697220 480 697460
rect 583520 697084 584960 697324
rect -960 684164 480 684404
rect 583520 683756 584960 683996
rect -960 671108 480 671348
rect 583520 670564 584960 670804
rect -960 658052 480 658292
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 583520 643908 584960 644148
rect -960 631940 480 632180
rect 583520 630716 584960 630956
rect -960 619020 480 619260
rect 583520 617388 584960 617628
rect -960 605964 480 606204
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 583520 590868 584960 591108
rect -960 579852 480 580092
rect 583520 577540 584960 577780
rect -960 566796 480 567036
rect 583520 564212 584960 564452
rect -960 553740 480 553980
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 583520 537692 584960 537932
rect -960 527764 480 528004
rect 583520 524364 584960 524604
rect -960 514708 480 514948
rect 583520 511172 584960 511412
rect -960 501652 480 501892
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 583520 484516 584960 484756
rect -960 475540 480 475780
rect 583520 471324 584960 471564
rect -960 462484 480 462724
rect 583520 457996 584960 458236
rect -960 449428 480 449668
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 583520 431476 584960 431716
rect -960 423452 480 423692
rect 583520 418148 584960 418388
rect -960 410396 480 410636
rect 583520 404820 584960 405060
rect -960 397340 480 397580
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 583520 378300 584960 378540
rect -960 371228 480 371468
rect 583520 364972 584960 365212
rect -960 358308 480 358548
rect 583520 351780 584960 352020
rect -960 345252 480 345492
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 583520 325124 584960 325364
rect -960 319140 480 319380
rect 583520 311932 584960 312172
rect -960 306084 480 306324
rect 583520 298604 584960 298844
rect -960 293028 480 293268
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 583520 272084 584960 272324
rect -960 267052 480 267292
rect 583520 258756 584960 258996
rect -960 253996 480 254236
rect 583520 245428 584960 245668
rect -960 240940 480 241180
rect 583520 232236 584960 232476
rect -960 227884 480 228124
rect 583520 218908 584960 219148
rect -960 214828 480 215068
rect 583520 205580 584960 205820
rect -960 201772 480 202012
rect 583520 192388 584960 192628
rect -960 188716 480 188956
rect 583520 179060 584960 179300
rect -960 175796 480 176036
rect 583520 165732 584960 165972
rect -960 162740 480 162980
rect 583520 152540 584960 152780
rect -960 149684 480 149924
rect 583520 139212 584960 139452
rect -960 136628 480 136868
rect 583520 125884 584960 126124
rect -960 123572 480 123812
rect 583520 112692 584960 112932
rect -960 110516 480 110756
rect 583520 99364 584960 99604
rect -960 97460 480 97700
rect 583520 86036 584960 86276
rect -960 84540 480 84780
rect 583520 72844 584960 73084
rect -960 71484 480 71724
rect 583520 59516 584960 59756
rect -960 58428 480 58668
rect 583520 46188 584960 46428
rect -960 45372 480 45612
rect 583520 32996 584960 33236
rect -960 32316 480 32556
rect 583520 19668 584960 19908
rect -960 19260 480 19500
rect -960 6340 480 6580
rect 583520 6476 584960 6716
<< obsm3 >>
rect 480 697540 583520 701793
rect 560 697404 583520 697540
rect 560 697140 583440 697404
rect 480 697004 583440 697140
rect 480 684484 583520 697004
rect 560 684084 583520 684484
rect 480 684076 583520 684084
rect 480 683676 583440 684076
rect 480 671428 583520 683676
rect 560 671028 583520 671428
rect 480 670884 583520 671028
rect 480 670484 583440 670884
rect 480 658372 583520 670484
rect 560 657972 583520 658372
rect 480 657556 583520 657972
rect 480 657156 583440 657556
rect 480 645316 583520 657156
rect 560 644916 583520 645316
rect 480 644228 583520 644916
rect 480 643828 583440 644228
rect 480 632260 583520 643828
rect 560 631860 583520 632260
rect 480 631036 583520 631860
rect 480 630636 583440 631036
rect 480 619340 583520 630636
rect 560 618940 583520 619340
rect 480 617708 583520 618940
rect 480 617308 583440 617708
rect 480 606284 583520 617308
rect 560 605884 583520 606284
rect 480 604380 583520 605884
rect 480 603980 583440 604380
rect 480 593228 583520 603980
rect 560 592828 583520 593228
rect 480 591188 583520 592828
rect 480 590788 583440 591188
rect 480 580172 583520 590788
rect 560 579772 583520 580172
rect 480 577860 583520 579772
rect 480 577460 583440 577860
rect 480 567116 583520 577460
rect 560 566716 583520 567116
rect 480 564532 583520 566716
rect 480 564132 583440 564532
rect 480 554060 583520 564132
rect 560 553660 583520 554060
rect 480 551340 583520 553660
rect 480 550940 583440 551340
rect 480 541004 583520 550940
rect 560 540604 583520 541004
rect 480 538012 583520 540604
rect 480 537612 583440 538012
rect 480 528084 583520 537612
rect 560 527684 583520 528084
rect 480 524684 583520 527684
rect 480 524284 583440 524684
rect 480 515028 583520 524284
rect 560 514628 583520 515028
rect 480 511492 583520 514628
rect 480 511092 583440 511492
rect 480 501972 583520 511092
rect 560 501572 583520 501972
rect 480 498164 583520 501572
rect 480 497764 583440 498164
rect 480 488916 583520 497764
rect 560 488516 583520 488916
rect 480 484836 583520 488516
rect 480 484436 583440 484836
rect 480 475860 583520 484436
rect 560 475460 583520 475860
rect 480 471644 583520 475460
rect 480 471244 583440 471644
rect 480 462804 583520 471244
rect 560 462404 583520 462804
rect 480 458316 583520 462404
rect 480 457916 583440 458316
rect 480 449748 583520 457916
rect 560 449348 583520 449748
rect 480 444988 583520 449348
rect 480 444588 583440 444988
rect 480 436828 583520 444588
rect 560 436428 583520 436828
rect 480 431796 583520 436428
rect 480 431396 583440 431796
rect 480 423772 583520 431396
rect 560 423372 583520 423772
rect 480 418468 583520 423372
rect 480 418068 583440 418468
rect 480 410716 583520 418068
rect 560 410316 583520 410716
rect 480 405140 583520 410316
rect 480 404740 583440 405140
rect 480 397660 583520 404740
rect 560 397260 583520 397660
rect 480 391948 583520 397260
rect 480 391548 583440 391948
rect 480 384604 583520 391548
rect 560 384204 583520 384604
rect 480 378620 583520 384204
rect 480 378220 583440 378620
rect 480 371548 583520 378220
rect 560 371148 583520 371548
rect 480 365292 583520 371148
rect 480 364892 583440 365292
rect 480 358628 583520 364892
rect 560 358228 583520 358628
rect 480 352100 583520 358228
rect 480 351700 583440 352100
rect 480 345572 583520 351700
rect 560 345172 583520 345572
rect 480 338772 583520 345172
rect 480 338372 583440 338772
rect 480 332516 583520 338372
rect 560 332116 583520 332516
rect 480 325444 583520 332116
rect 480 325044 583440 325444
rect 480 319460 583520 325044
rect 560 319060 583520 319460
rect 480 312252 583520 319060
rect 480 311852 583440 312252
rect 480 306404 583520 311852
rect 560 306004 583520 306404
rect 480 298924 583520 306004
rect 480 298524 583440 298924
rect 480 293348 583520 298524
rect 560 292948 583520 293348
rect 480 285596 583520 292948
rect 480 285196 583440 285596
rect 480 280292 583520 285196
rect 560 279892 583520 280292
rect 480 272404 583520 279892
rect 480 272004 583440 272404
rect 480 267372 583520 272004
rect 560 266972 583520 267372
rect 480 259076 583520 266972
rect 480 258676 583440 259076
rect 480 254316 583520 258676
rect 560 253916 583520 254316
rect 480 245748 583520 253916
rect 480 245348 583440 245748
rect 480 241260 583520 245348
rect 560 240860 583520 241260
rect 480 232556 583520 240860
rect 480 232156 583440 232556
rect 480 228204 583520 232156
rect 560 227804 583520 228204
rect 480 219228 583520 227804
rect 480 218828 583440 219228
rect 480 215148 583520 218828
rect 560 214748 583520 215148
rect 480 205900 583520 214748
rect 480 205500 583440 205900
rect 480 202092 583520 205500
rect 560 201692 583520 202092
rect 480 192708 583520 201692
rect 480 192308 583440 192708
rect 480 189036 583520 192308
rect 560 188636 583520 189036
rect 480 179380 583520 188636
rect 480 178980 583440 179380
rect 480 176116 583520 178980
rect 560 175716 583520 176116
rect 480 166052 583520 175716
rect 480 165652 583440 166052
rect 480 163060 583520 165652
rect 560 162660 583520 163060
rect 480 152860 583520 162660
rect 480 152460 583440 152860
rect 480 150004 583520 152460
rect 560 149604 583520 150004
rect 480 139532 583520 149604
rect 480 139132 583440 139532
rect 480 136948 583520 139132
rect 560 136548 583520 136948
rect 480 126204 583520 136548
rect 480 125804 583440 126204
rect 480 123892 583520 125804
rect 560 123492 583520 123892
rect 480 113012 583520 123492
rect 480 112612 583440 113012
rect 480 110836 583520 112612
rect 560 110436 583520 110836
rect 480 99684 583520 110436
rect 480 99284 583440 99684
rect 480 97780 583520 99284
rect 560 97380 583520 97780
rect 480 86356 583520 97380
rect 480 85956 583440 86356
rect 480 84860 583520 85956
rect 560 84460 583520 84860
rect 480 73164 583520 84460
rect 480 72764 583440 73164
rect 480 71804 583520 72764
rect 560 71404 583520 71804
rect 480 59836 583520 71404
rect 480 59436 583440 59836
rect 480 58748 583520 59436
rect 560 58348 583520 58748
rect 480 46508 583520 58348
rect 480 46108 583440 46508
rect 480 45692 583520 46108
rect 560 45292 583520 45692
rect 480 33316 583520 45292
rect 480 32916 583440 33316
rect 480 32636 583520 32916
rect 560 32236 583520 32636
rect 480 19988 583520 32236
rect 480 19588 583440 19988
rect 480 19580 583520 19588
rect 560 19180 583520 19580
rect 480 6796 583520 19180
rect 480 6660 583440 6796
rect 560 6396 583440 6660
rect 560 6260 583520 6396
rect 480 2143 583520 6260
<< metal4 >>
rect 1794 2128 2414 701808
rect 5514 2128 6134 701808
rect 9234 2128 9854 701808
rect 12954 2128 13574 701808
rect 16674 2128 17294 701808
rect 20394 2128 21014 701808
rect 24114 2128 24734 701808
rect 27834 2128 28454 701808
rect 37794 670412 38414 701808
rect 41514 670412 42134 701808
rect 73794 670412 74414 701808
rect 77514 670412 78134 701808
rect 109794 670412 110414 701808
rect 113514 670412 114134 701808
rect 37794 546808 38414 577112
rect 41514 546808 42134 577112
rect 73794 546808 74414 577112
rect 77514 546808 78134 577112
rect 109794 546808 110414 577112
rect 113514 546808 114134 577112
rect 135834 546808 136454 701808
rect 37794 431364 38414 462212
rect 41514 431364 42134 462212
rect 73794 431364 74414 462088
rect 77514 431488 78134 462088
rect 109794 431488 110414 462212
rect 113514 431364 114134 462212
rect 145794 431364 146414 701808
rect 149514 431364 150134 701808
rect 153234 431364 153854 701808
rect 156954 431364 157574 701808
rect 160674 431364 161294 701808
rect 164394 431364 165014 701808
rect 168114 431364 168734 701808
rect 171834 431364 172454 701808
rect 181794 431364 182414 701808
rect 37794 201136 38414 293048
rect 41514 201136 42134 293048
rect 45234 201136 45854 293048
rect 48954 201136 49574 293048
rect 52674 201136 53294 293048
rect 56394 201136 57014 292924
rect 60114 201136 60734 292924
rect 63834 201136 64454 292924
rect 73794 201136 74414 292924
rect 77514 201260 78134 292924
rect 81234 201136 81854 293048
rect 84954 201260 85574 292924
rect 88674 201136 89294 292924
rect 92394 201260 93014 292924
rect 96114 201136 96734 292924
rect 99834 201260 100454 292924
rect 109794 201260 110414 292924
rect 113514 201136 114134 293048
rect 117234 201260 117854 292924
rect 120954 201136 121574 293048
rect 124674 201260 125294 292924
rect 128394 201136 129014 293048
rect 132114 201260 132734 292924
rect 135834 201136 136454 293048
rect 145794 201136 146414 293048
rect 149514 201136 150134 293048
rect 153234 201136 153854 293048
rect 156954 201136 157574 293048
rect 160674 201260 161294 293048
rect 164394 201136 165014 293048
rect 168114 201136 168734 293048
rect 171834 201136 172454 293048
rect 37794 82020 38414 113548
rect 41514 82020 42134 113548
rect 73794 82020 74414 113424
rect 77514 82020 78134 113424
rect 109794 82020 110414 113548
rect 113514 82020 114134 113548
rect 37794 2128 38414 33464
rect 41514 2128 42134 33464
rect 73794 2128 74414 33340
rect 77514 2128 78134 33340
rect 109794 2128 110414 33464
rect 113514 2128 114134 33464
rect 145794 2128 146414 113548
rect 149514 2128 150134 113548
rect 153234 2128 153854 113548
rect 156954 2128 157574 113548
rect 160674 2128 161294 113548
rect 164394 2128 165014 113548
rect 168114 2128 168734 113548
rect 171834 2128 172454 113548
rect 181794 2128 182414 293048
rect 185514 2128 186134 701808
rect 189234 2128 189854 701808
rect 192954 2128 193574 701808
rect 196674 2128 197294 701808
rect 200394 2128 201014 701808
rect 204114 2128 204734 701808
rect 207834 2128 208454 701808
rect 217794 2128 218414 701808
rect 221514 2128 222134 701808
rect 225234 2128 225854 701808
rect 228954 2128 229574 701808
rect 232674 2128 233294 701808
rect 236394 2128 237014 701808
rect 240114 2128 240734 701808
rect 243834 2128 244454 701808
rect 253794 2128 254414 701808
rect 257514 2128 258134 701808
rect 261234 2128 261854 701808
rect 264954 2128 265574 701808
rect 268674 2128 269294 701808
rect 272394 2128 273014 701808
rect 276114 2128 276734 701808
rect 279834 2128 280454 701808
rect 289794 2128 290414 701808
rect 293514 2128 294134 701808
rect 297234 2128 297854 701808
rect 300954 2128 301574 701808
rect 304674 2128 305294 701808
rect 308394 2128 309014 701808
rect 312114 2128 312734 701808
rect 315834 2128 316454 701808
rect 325794 122660 326414 701808
rect 329514 122660 330134 701808
rect 333234 122660 333854 701808
rect 336954 122660 337574 701808
rect 361794 672944 362414 701808
rect 365514 672944 366134 701808
rect 397794 672944 398414 701808
rect 401514 672944 402134 701808
rect 433794 672944 434414 701808
rect 437514 672944 438134 701808
rect 340674 548516 341294 603852
rect 344394 548516 345014 603852
rect 348114 548516 348734 603852
rect 361794 548516 362414 603728
rect 365514 548516 366134 603728
rect 369234 548516 369854 603728
rect 372954 548640 373574 603852
rect 376674 548516 377294 603852
rect 380394 548640 381014 603728
rect 384114 548516 384734 603728
rect 397794 548640 398414 603728
rect 401514 548516 402134 603728
rect 405234 548640 405854 603728
rect 408954 548516 409574 603852
rect 412674 548640 413294 603852
rect 416394 548516 417014 603852
rect 420114 548640 420734 603852
rect 433794 548516 434414 603852
rect 437514 548640 438134 603852
rect 441234 548516 441854 701808
rect 444954 548640 445574 701808
rect 448674 548516 449294 701808
rect 452394 548516 453014 701808
rect 456114 548516 456734 701808
rect 459834 548516 460454 701808
rect 469794 548516 470414 701808
rect 473514 548640 474134 701808
rect 477234 548516 477854 701808
rect 480954 548516 481574 701808
rect 361794 368088 362414 410076
rect 365514 368088 366134 410076
rect 369234 368088 369854 410076
rect 372954 368088 373574 410076
rect 397794 368088 398414 410076
rect 401514 368088 402134 410200
rect 405234 368088 405854 410076
rect 408954 368088 409574 410200
rect 433794 368088 434414 410200
rect 437514 368088 438134 410076
rect 351834 244852 352454 298996
rect 361794 244852 362414 298872
rect 365514 244852 366134 298872
rect 369234 244976 369854 298872
rect 387834 244852 388454 298872
rect 397794 244852 398414 298872
rect 401514 244852 402134 298872
rect 405234 244852 405854 298872
rect 423834 244852 424454 298872
rect 433794 244852 434414 298996
rect 437514 244852 438134 298996
rect 441234 244852 441854 410200
rect 444954 244852 445574 410076
rect 448674 244852 449294 410200
rect 452394 244852 453014 410200
rect 456114 244852 456734 410200
rect 459834 244852 460454 410200
rect 469794 244852 470414 410200
rect 473514 244852 474134 410200
rect 477234 244852 477854 410200
rect 361794 122784 362414 157140
rect 365514 122784 366134 157140
rect 397794 122660 398414 157140
rect 401514 122784 402134 157264
rect 325794 2128 326414 38064
rect 329514 2128 330134 38064
rect 361794 2128 362414 37940
rect 365514 2128 366134 37940
rect 397794 2128 398414 38064
rect 401514 2128 402134 38064
rect 423834 2128 424454 157264
rect 433794 2128 434414 157264
rect 437514 2128 438134 157264
rect 441234 2128 441854 157264
rect 444954 2128 445574 157264
rect 448674 2128 449294 157264
rect 452394 2128 453014 157264
rect 469794 122660 470414 157264
rect 473514 122660 474134 157264
rect 480954 122660 481574 410200
rect 484674 122784 485294 701808
rect 488394 122660 489014 701808
rect 492114 122660 492734 701808
rect 495834 122660 496454 701808
rect 505794 655298 506414 701808
rect 505794 122660 506414 603728
rect 509514 122660 510134 701808
rect 513234 122660 513854 701808
rect 516954 122660 517574 701808
rect 520674 122660 521294 701808
rect 524394 122660 525014 701808
rect 528114 122660 528734 701808
rect 531834 122660 532454 701808
rect 541794 122660 542414 701808
rect 545514 122660 546134 701808
rect 549234 122660 549854 701808
rect 552954 122660 553574 701808
rect 469794 2128 470414 38064
rect 473514 2128 474134 37940
rect 505794 2128 506414 37940
rect 509514 2128 510134 38064
rect 541794 2128 542414 38064
rect 545514 2128 546134 38064
rect 556674 2128 557294 701808
rect 560394 2128 561014 701808
rect 564114 2128 564734 701808
rect 567834 2128 568454 701808
rect 577794 2128 578414 701808
rect 581514 2128 582134 701808
<< obsm4 >>
rect 35755 670332 37714 671125
rect 38494 670332 41434 671125
rect 42214 670332 73714 671125
rect 74494 670332 77434 671125
rect 78214 670332 109714 671125
rect 110494 670332 113434 671125
rect 114214 670332 135754 671125
rect 35755 577192 135754 670332
rect 35755 546728 37714 577192
rect 38494 546728 41434 577192
rect 42214 546728 73714 577192
rect 74494 546728 77434 577192
rect 78214 546728 109714 577192
rect 110494 546728 113434 577192
rect 114214 546728 135754 577192
rect 136534 546728 145714 671125
rect 35755 462292 145714 546728
rect 35755 431284 37714 462292
rect 38494 431284 41434 462292
rect 42214 462168 109714 462292
rect 42214 431284 73714 462168
rect 74494 431408 77434 462168
rect 78214 431408 109714 462168
rect 110494 431408 113434 462292
rect 74494 431284 113434 431408
rect 114214 431284 145714 462292
rect 146494 431284 149434 671125
rect 150214 431284 153154 671125
rect 153934 431284 156874 671125
rect 157654 431284 160594 671125
rect 161374 431284 164314 671125
rect 165094 431284 168034 671125
rect 168814 431284 171754 671125
rect 172534 431284 181714 671125
rect 182494 431284 185434 671125
rect 35755 293128 185434 431284
rect 35755 201056 37714 293128
rect 38494 201056 41434 293128
rect 42214 201056 45154 293128
rect 45934 201056 48874 293128
rect 49654 201056 52594 293128
rect 53374 293004 81154 293128
rect 53374 201056 56314 293004
rect 57094 201056 60034 293004
rect 60814 201056 63754 293004
rect 64534 201056 73714 293004
rect 74494 201180 77434 293004
rect 78214 201180 81154 293004
rect 74494 201056 81154 201180
rect 81934 293004 113434 293128
rect 81934 201180 84874 293004
rect 85654 201180 88594 293004
rect 81934 201056 88594 201180
rect 89374 201180 92314 293004
rect 93094 201180 96034 293004
rect 89374 201056 96034 201180
rect 96814 201180 99754 293004
rect 100534 201180 109714 293004
rect 110494 201180 113434 293004
rect 96814 201056 113434 201180
rect 114214 293004 120874 293128
rect 114214 201180 117154 293004
rect 117934 201180 120874 293004
rect 114214 201056 120874 201180
rect 121654 293004 128314 293128
rect 121654 201180 124594 293004
rect 125374 201180 128314 293004
rect 121654 201056 128314 201180
rect 129094 293004 135754 293128
rect 129094 201180 132034 293004
rect 132814 201180 135754 293004
rect 129094 201056 135754 201180
rect 136534 201056 145714 293128
rect 146494 201056 149434 293128
rect 150214 201056 153154 293128
rect 153934 201056 156874 293128
rect 157654 201180 160594 293128
rect 161374 201180 164314 293128
rect 157654 201056 164314 201180
rect 165094 201056 168034 293128
rect 168814 201056 171754 293128
rect 172534 201056 181714 293128
rect 35755 113628 181714 201056
rect 35755 81940 37714 113628
rect 38494 81940 41434 113628
rect 42214 113504 109714 113628
rect 42214 81940 73714 113504
rect 74494 81940 77434 113504
rect 78214 81940 109714 113504
rect 110494 81940 113434 113628
rect 114214 81940 145714 113628
rect 35755 33544 145714 81940
rect 35755 17171 37714 33544
rect 38494 17171 41434 33544
rect 42214 33420 109714 33544
rect 42214 17171 73714 33420
rect 74494 17171 77434 33420
rect 78214 17171 109714 33420
rect 110494 17171 113434 33544
rect 114214 17171 145714 33544
rect 146494 17171 149434 113628
rect 150214 17171 153154 113628
rect 153934 17171 156874 113628
rect 157654 17171 160594 113628
rect 161374 17171 164314 113628
rect 165094 17171 168034 113628
rect 168814 17171 171754 113628
rect 172534 17171 181714 113628
rect 182494 17171 185434 293128
rect 186214 17171 189154 671125
rect 189934 17171 192874 671125
rect 193654 17171 196594 671125
rect 197374 17171 200314 671125
rect 201094 17171 204034 671125
rect 204814 17171 207754 671125
rect 208534 17171 217714 671125
rect 218494 17171 221434 671125
rect 222214 17171 225154 671125
rect 225934 17171 228874 671125
rect 229654 17171 232594 671125
rect 233374 17171 236314 671125
rect 237094 17171 240034 671125
rect 240814 17171 243754 671125
rect 244534 17171 253714 671125
rect 254494 17171 257434 671125
rect 258214 17171 261154 671125
rect 261934 17171 264874 671125
rect 265654 17171 268594 671125
rect 269374 17171 272314 671125
rect 273094 17171 276034 671125
rect 276814 17171 279754 671125
rect 280534 17171 289714 671125
rect 290494 17171 293434 671125
rect 294214 17171 297154 671125
rect 297934 17171 300874 671125
rect 301654 17171 304594 671125
rect 305374 17171 308314 671125
rect 309094 17171 312034 671125
rect 312814 17171 315754 671125
rect 316534 122580 325714 671125
rect 326494 122580 329434 671125
rect 330214 122580 333154 671125
rect 333934 122580 336874 671125
rect 337654 603932 441154 671125
rect 337654 548436 340594 603932
rect 341374 548436 344314 603932
rect 345094 548436 348034 603932
rect 348814 603808 372874 603932
rect 348814 548436 361714 603808
rect 362494 548436 365434 603808
rect 366214 548436 369154 603808
rect 369934 548560 372874 603808
rect 373654 548560 376594 603932
rect 369934 548436 376594 548560
rect 377374 603808 408874 603932
rect 377374 548560 380314 603808
rect 381094 548560 384034 603808
rect 377374 548436 384034 548560
rect 384814 548560 397714 603808
rect 398494 548560 401434 603808
rect 384814 548436 401434 548560
rect 402214 548560 405154 603808
rect 405934 548560 408874 603808
rect 402214 548436 408874 548560
rect 409654 548560 412594 603932
rect 413374 548560 416314 603932
rect 409654 548436 416314 548560
rect 417094 548560 420034 603932
rect 420814 548560 433714 603932
rect 417094 548436 433714 548560
rect 434494 548560 437434 603932
rect 438214 548560 441154 603932
rect 434494 548436 441154 548560
rect 441934 548560 444874 671125
rect 445654 548560 448594 671125
rect 441934 548436 448594 548560
rect 449374 548436 452314 671125
rect 453094 548436 456034 671125
rect 456814 548436 459754 671125
rect 460534 548436 469714 671125
rect 470494 548560 473434 671125
rect 474214 548560 477154 671125
rect 470494 548436 477154 548560
rect 477934 548436 480874 671125
rect 481654 548436 484594 671125
rect 337654 410280 484594 548436
rect 337654 410156 401434 410280
rect 337654 368008 361714 410156
rect 362494 368008 365434 410156
rect 366214 368008 369154 410156
rect 369934 368008 372874 410156
rect 373654 368008 397714 410156
rect 398494 368008 401434 410156
rect 402214 410156 408874 410280
rect 402214 368008 405154 410156
rect 405934 368008 408874 410156
rect 409654 368008 433714 410280
rect 434494 410156 441154 410280
rect 434494 368008 437434 410156
rect 438214 368008 441154 410156
rect 337654 299076 441154 368008
rect 337654 244772 351754 299076
rect 352534 298952 433714 299076
rect 352534 244772 361714 298952
rect 362494 244772 365434 298952
rect 366214 244896 369154 298952
rect 369934 244896 387754 298952
rect 366214 244772 387754 244896
rect 388534 244772 397714 298952
rect 398494 244772 401434 298952
rect 402214 244772 405154 298952
rect 405934 244772 423754 298952
rect 424534 244772 433714 298952
rect 434494 244772 437434 299076
rect 438214 244772 441154 299076
rect 441934 410156 448594 410280
rect 441934 244772 444874 410156
rect 445654 244772 448594 410156
rect 449374 244772 452314 410280
rect 453094 244772 456034 410280
rect 456814 244772 459754 410280
rect 460534 244772 469714 410280
rect 470494 244772 473434 410280
rect 474214 244772 477154 410280
rect 477934 244772 480874 410280
rect 337654 157344 480874 244772
rect 337654 157220 401434 157344
rect 337654 122704 361714 157220
rect 362494 122704 365434 157220
rect 366214 122704 397714 157220
rect 337654 122580 397714 122704
rect 398494 122704 401434 157220
rect 402214 122704 423754 157344
rect 398494 122580 423754 122704
rect 316534 38144 423754 122580
rect 316534 17171 325714 38144
rect 326494 17171 329434 38144
rect 330214 38020 397714 38144
rect 330214 17171 361714 38020
rect 362494 17171 365434 38020
rect 366214 17171 397714 38020
rect 398494 17171 401434 38144
rect 402214 17171 423754 38144
rect 424534 17171 433714 157344
rect 434494 17171 437434 157344
rect 438214 17171 441154 157344
rect 441934 17171 444874 157344
rect 445654 17171 448594 157344
rect 449374 17171 452314 157344
rect 453094 122580 469714 157344
rect 470494 122580 473434 157344
rect 474214 122580 480874 157344
rect 481654 122704 484594 410280
rect 485374 122704 488314 671125
rect 481654 122580 488314 122704
rect 489094 122580 492034 671125
rect 492814 122580 495754 671125
rect 496534 655218 505714 671125
rect 506494 655218 509434 671125
rect 496534 603808 509434 655218
rect 496534 122580 505714 603808
rect 506494 122580 509434 603808
rect 510214 122580 513154 671125
rect 513934 122580 516874 671125
rect 517654 122580 520594 671125
rect 521374 122580 524314 671125
rect 525094 122580 528034 671125
rect 528814 122580 531754 671125
rect 532534 122580 541714 671125
rect 542494 122580 545434 671125
rect 546214 122580 549154 671125
rect 549934 122580 552874 671125
rect 553654 122580 554632 671125
rect 453094 38144 554632 122580
rect 453094 17171 469714 38144
rect 470494 38020 509434 38144
rect 470494 17171 473434 38020
rect 474214 17171 505714 38020
rect 506494 17171 509434 38020
rect 510214 17171 541714 38144
rect 542494 17171 545434 38144
rect 546214 17171 554632 38144
<< metal5 >>
rect 1056 698026 582868 698646
rect 1056 694306 582868 694926
rect 1056 690586 582868 691206
rect 1056 686866 582868 687486
rect 1056 676906 582868 677526
rect 1056 673186 582868 673806
rect 1056 669466 582868 670086
rect 1056 665746 582868 666366
rect 1056 662026 582868 662646
rect 1056 658306 582868 658926
rect 1056 654586 582868 655206
rect 1056 650866 582868 651486
rect 1056 640906 582868 641526
rect 1056 637186 582868 637806
rect 1056 633466 582868 634086
rect 1056 629746 582868 630366
rect 1056 626026 582868 626646
rect 1056 622306 582868 622926
rect 1056 618586 582868 619206
rect 1056 614866 582868 615486
rect 1056 604906 582868 605526
rect 1056 601186 582868 601806
rect 1056 597466 582868 598086
rect 1056 593746 582868 594366
rect 1056 590026 582868 590646
rect 1056 586306 582868 586926
rect 1056 582586 582868 583206
rect 1056 578866 582868 579486
rect 1056 568906 582868 569526
rect 1056 565186 582868 565806
rect 1056 561466 582868 562086
rect 1056 557746 582868 558366
rect 1056 554026 582868 554646
rect 1056 550306 582868 550926
rect 1794 548110 146414 548730
rect 1056 546586 582868 547206
rect 1056 542866 582868 543486
rect 1056 532906 582868 533526
rect 1056 529186 582868 529806
rect 1056 525466 582868 526086
rect 1056 521746 582868 522366
rect 1056 518026 582868 518646
rect 1056 514306 582868 514926
rect 1056 510586 582868 511206
rect 1056 506866 582868 507486
rect 1056 496906 582868 497526
rect 1056 493186 582868 493806
rect 1056 489466 582868 490086
rect 1056 485746 582868 486366
rect 1056 482026 582868 482646
rect 1056 478306 582868 478926
rect 1056 474586 582868 475206
rect 1056 470866 582868 471486
rect 1056 460906 582868 461526
rect 1056 457186 582868 457806
rect 1056 453466 582868 454086
rect 1056 449746 582868 450366
rect 1056 446026 582868 446646
rect 1056 442306 582868 442926
rect 1056 438586 582868 439206
rect 1056 434866 582868 435486
rect 1056 424906 582868 425526
rect 1056 421186 582868 421806
rect 1056 417466 582868 418086
rect 1056 413746 582868 414366
rect 1056 410026 582868 410646
rect 1056 406306 582868 406926
rect 1056 402586 582868 403206
rect 1056 398866 582868 399486
rect 1056 388906 582868 389526
rect 1056 385186 582868 385806
rect 1056 381466 582868 382086
rect 1056 377746 582868 378366
rect 1056 374026 582868 374646
rect 1056 370306 582868 370926
rect 1056 366586 582868 367206
rect 1056 362866 582868 363486
rect 1056 352906 582868 353526
rect 1056 349186 582868 349806
rect 1056 345466 582868 346086
rect 1056 341746 582868 342366
rect 1056 338026 582868 338646
rect 1056 334306 582868 334926
rect 1056 330586 582868 331206
rect 1056 326866 582868 327486
rect 1056 316906 582868 317526
rect 1056 313186 582868 313806
rect 1056 309466 582868 310086
rect 1056 305746 582868 306366
rect 1056 302026 582868 302646
rect 1056 298306 582868 298926
rect 1056 294586 582868 295206
rect 1056 290866 582868 291486
rect 1056 280906 582868 281526
rect 1056 277186 582868 277806
rect 1056 273466 582868 274086
rect 1056 269746 582868 270366
rect 1056 266026 582868 266646
rect 1056 262306 582868 262926
rect 1056 258586 582868 259206
rect 1056 254866 582868 255486
rect 1056 244906 582868 245526
rect 1056 241186 582868 241806
rect 1056 237466 582868 238086
rect 1056 233746 582868 234366
rect 1056 230026 582868 230646
rect 1056 226306 582868 226926
rect 1056 222586 582868 223206
rect 1056 218866 582868 219486
rect 1056 208906 582868 209526
rect 1056 205186 582868 205806
rect 1056 201466 582868 202086
rect 1056 197746 582868 198366
rect 1056 194026 582868 194646
rect 1056 190306 582868 190926
rect 1056 186586 582868 187206
rect 1056 182866 582868 183486
rect 1056 172906 582868 173526
rect 1056 169186 582868 169806
rect 1056 165466 582868 166086
rect 1056 161746 582868 162366
rect 1056 158026 582868 158646
rect 1056 154306 582868 154926
rect 1056 150586 582868 151206
rect 1056 146866 582868 147486
rect 1056 136906 582868 137526
rect 1056 133186 582868 133806
rect 1056 129466 582868 130086
rect 1056 125746 582868 126366
rect 1056 122026 582868 122646
rect 1056 118306 582868 118926
rect 1056 114586 582868 115206
rect 1056 110866 582868 111486
rect 1056 100906 582868 101526
rect 1056 97186 582868 97806
rect 1056 93466 582868 94086
rect 1056 89746 582868 90366
rect 1056 86026 582868 86646
rect 5514 83670 150134 84290
rect 1056 82306 582868 82926
rect 1056 78586 582868 79206
rect 1056 74866 582868 75486
rect 1056 64906 582868 65526
rect 1056 61186 582868 61806
rect 1056 57466 582868 58086
rect 1056 53746 582868 54366
rect 1056 50026 582868 50646
rect 1056 46306 582868 46926
rect 1056 42586 582868 43206
rect 1056 38866 582868 39486
rect 1056 28906 582868 29526
rect 1056 25186 582868 25806
rect 1056 21466 582868 22086
rect 1056 17746 582868 18366
rect 1056 14026 582868 14646
rect 1056 10306 582868 10926
rect 1056 6586 582868 7206
rect 1056 2866 582868 3486
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 1 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 2 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 3 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 4 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 5 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 6 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 7 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 8 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 9 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 10 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 11 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 12 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 13 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 14 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 15 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 16 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 17 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 18 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 19 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 20 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 26 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 27 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 28 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 29 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 30 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 32 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 33 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 34 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 35 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 36 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 37 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 38 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 39 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 40 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 41 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 42 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 43 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 44 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 45 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 46 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 47 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 48 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 49 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 50 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 51 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 52 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 53 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 54 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 55 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 56 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 57 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 58 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 59 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 60 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 61 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 62 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 63 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 64 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 65 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 66 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 67 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 68 nsew signal output
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 69 nsew signal output
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 70 nsew signal output
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 71 nsew signal output
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 72 nsew signal output
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 73 nsew signal output
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 74 nsew signal output
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 75 nsew signal output
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 76 nsew signal output
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 77 nsew signal output
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 78 nsew signal output
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 79 nsew signal output
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 80 nsew signal output
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 81 nsew signal output
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 82 nsew signal output
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 83 nsew signal output
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 84 nsew signal output
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 85 nsew signal output
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 86 nsew signal output
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 87 nsew signal output
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 88 nsew signal output
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 89 nsew signal output
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 90 nsew signal output
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 91 nsew signal output
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 92 nsew signal output
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 93 nsew signal output
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 94 nsew signal output
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 95 nsew signal output
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 96 nsew signal output
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 97 nsew signal output
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 98 nsew signal output
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 99 nsew signal output
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 100 nsew signal output
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 101 nsew signal output
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 102 nsew signal output
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 103 nsew signal output
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 104 nsew signal output
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 105 nsew signal output
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 106 nsew signal output
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 107 nsew signal output
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 108 nsew signal output
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 109 nsew signal output
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 110 nsew signal output
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 111 nsew signal output
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 112 nsew signal output
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 113 nsew signal output
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 114 nsew signal output
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 115 nsew signal output
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 116 nsew signal output
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 117 nsew signal output
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 118 nsew signal output
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 119 nsew signal output
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 120 nsew signal output
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 121 nsew signal output
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 122 nsew signal output
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 123 nsew signal output
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 124 nsew signal output
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 125 nsew signal output
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 126 nsew signal output
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 127 nsew signal output
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 128 nsew signal output
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 129 nsew signal output
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 130 nsew signal output
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 131 nsew signal output
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 132 nsew signal output
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 133 nsew signal output
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 134 nsew signal output
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 135 nsew signal output
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 136 nsew signal output
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 137 nsew signal output
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 138 nsew signal output
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 139 nsew signal output
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 140 nsew signal output
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 141 nsew signal output
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 142 nsew signal output
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 143 nsew signal output
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 144 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 145 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 146 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 147 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 148 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 149 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 150 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 151 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 152 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 153 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 154 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 155 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 156 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 157 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 158 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 159 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 160 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 161 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 162 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 163 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 164 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 165 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 166 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 167 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 168 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 169 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 170 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 171 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 172 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 173 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 174 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 175 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 176 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 177 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 178 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 179 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 180 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 181 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 182 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 183 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 184 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 185 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 186 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 187 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 188 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 189 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 190 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 191 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 192 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 193 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 194 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 195 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 196 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 197 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 198 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 199 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 200 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 201 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 202 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 203 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 204 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 205 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 206 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 207 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 208 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 209 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 210 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 211 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 212 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 213 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 214 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 215 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 216 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 217 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 218 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 219 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 220 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 221 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 222 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 223 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 224 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 225 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 226 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 227 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 228 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 229 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 230 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 231 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 232 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 233 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 234 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 235 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 236 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 237 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 238 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 239 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 240 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 241 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 242 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 243 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 244 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 245 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 246 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 247 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 248 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 249 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 250 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 251 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 252 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 253 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 254 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 255 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 256 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 257 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 258 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 259 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 260 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 261 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 262 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 263 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 264 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 265 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 266 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 267 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 268 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 269 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 270 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 271 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 272 nsew signal output
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 273 nsew signal output
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 274 nsew signal output
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 275 nsew signal output
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 276 nsew signal output
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 277 nsew signal output
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 278 nsew signal output
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 279 nsew signal output
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 280 nsew signal output
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 281 nsew signal output
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 282 nsew signal output
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 283 nsew signal output
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 284 nsew signal output
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 285 nsew signal output
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 286 nsew signal output
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 287 nsew signal output
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 288 nsew signal output
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 289 nsew signal output
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 290 nsew signal output
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 291 nsew signal output
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 292 nsew signal output
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 293 nsew signal output
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 294 nsew signal output
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 295 nsew signal output
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 296 nsew signal output
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 297 nsew signal output
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 298 nsew signal output
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 299 nsew signal output
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 300 nsew signal output
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 301 nsew signal output
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 302 nsew signal output
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 303 nsew signal output
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 304 nsew signal output
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 305 nsew signal output
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 306 nsew signal output
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 307 nsew signal output
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 308 nsew signal output
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 309 nsew signal output
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 310 nsew signal output
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 311 nsew signal output
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 312 nsew signal output
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 313 nsew signal output
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 314 nsew signal output
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 315 nsew signal output
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 316 nsew signal output
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 317 nsew signal output
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 318 nsew signal output
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 319 nsew signal output
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 320 nsew signal output
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 321 nsew signal output
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 322 nsew signal output
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 323 nsew signal output
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 324 nsew signal output
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 325 nsew signal output
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 326 nsew signal output
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 327 nsew signal output
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 328 nsew signal output
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 329 nsew signal output
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 330 nsew signal output
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 331 nsew signal output
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 332 nsew signal output
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 333 nsew signal output
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 334 nsew signal output
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 335 nsew signal output
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 336 nsew signal output
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 337 nsew signal output
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 338 nsew signal output
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 339 nsew signal output
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 340 nsew signal output
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 341 nsew signal output
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 342 nsew signal output
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 343 nsew signal output
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 344 nsew signal output
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 345 nsew signal output
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 346 nsew signal output
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 347 nsew signal output
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 348 nsew signal output
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 349 nsew signal output
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 350 nsew signal output
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 351 nsew signal output
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 352 nsew signal output
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 353 nsew signal output
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 354 nsew signal output
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 355 nsew signal output
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 356 nsew signal output
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 357 nsew signal output
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 358 nsew signal output
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 359 nsew signal output
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 360 nsew signal output
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 361 nsew signal output
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 362 nsew signal output
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 363 nsew signal output
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 364 nsew signal output
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 365 nsew signal output
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 366 nsew signal output
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 367 nsew signal output
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 368 nsew signal output
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 369 nsew signal output
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 370 nsew signal output
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 371 nsew signal output
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 372 nsew signal output
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 373 nsew signal output
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 374 nsew signal output
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 375 nsew signal output
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 376 nsew signal output
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 377 nsew signal output
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 378 nsew signal output
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 379 nsew signal output
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 380 nsew signal output
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 381 nsew signal output
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 382 nsew signal output
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 383 nsew signal output
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 384 nsew signal output
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 385 nsew signal output
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 386 nsew signal output
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 387 nsew signal output
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 388 nsew signal output
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 389 nsew signal output
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 390 nsew signal output
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 391 nsew signal output
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 392 nsew signal output
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 393 nsew signal output
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 394 nsew signal output
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 395 nsew signal output
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 396 nsew signal output
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 397 nsew signal output
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 398 nsew signal output
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 399 nsew signal output
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 400 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 401 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 402 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 403 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 404 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 405 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 406 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 407 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 408 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 409 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 410 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 411 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 412 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 413 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 414 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 415 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 416 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 417 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 418 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 419 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 420 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 421 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 422 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 423 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 424 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 425 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 426 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 427 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 428 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 429 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 430 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 431 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 432 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 433 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 434 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 435 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 436 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 437 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 438 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 439 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 440 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 441 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 442 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 443 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 444 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 445 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 446 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 447 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 448 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 449 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 450 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 451 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 452 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 453 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 454 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 455 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 456 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 457 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 458 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 459 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 460 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 461 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 462 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 463 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 464 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 465 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 466 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 467 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 468 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 469 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 470 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 471 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 472 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 473 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 474 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 475 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 476 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 477 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 478 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 479 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 480 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 481 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 482 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 483 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 484 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 485 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 486 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 487 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 488 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 489 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 490 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 491 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 492 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 493 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 494 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 495 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 496 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 497 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 498 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 499 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 500 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 501 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 502 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 503 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 504 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 505 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 506 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 507 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 508 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 509 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 510 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 511 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 512 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 513 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 514 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 515 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 516 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 517 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 518 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 519 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 520 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 521 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 522 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 523 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 524 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 525 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 526 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 527 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 528 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 529 nsew signal output
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 530 nsew signal output
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 531 nsew signal output
rlabel metal4 s 1794 2128 2414 701808 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 37794 2128 38414 33464 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 37794 82020 38414 113548 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 37794 201136 38414 293048 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 37794 431364 38414 462212 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 37794 546808 38414 577112 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 37794 670412 38414 701808 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 73794 2128 74414 33340 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 73794 82020 74414 113424 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 73794 201136 74414 292924 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 73794 431364 74414 462088 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 73794 546808 74414 577112 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 73794 670412 74414 701808 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 109794 2128 110414 33464 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 109794 82020 110414 113548 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 109794 201260 110414 292924 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 109794 431488 110414 462212 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 109794 546808 110414 577112 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 109794 670412 110414 701808 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 145794 2128 146414 113548 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 145794 201136 146414 293048 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 145794 431364 146414 701808 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 181794 2128 182414 293048 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 181794 431364 182414 701808 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 217794 2128 218414 701808 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 253794 2128 254414 701808 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 289794 2128 290414 701808 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 325794 2128 326414 38064 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 325794 122660 326414 701808 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 361794 2128 362414 37940 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 361794 122784 362414 157140 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 361794 244852 362414 298872 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 361794 368088 362414 410076 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 361794 548516 362414 603728 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 361794 672944 362414 701808 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 397794 2128 398414 38064 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 397794 122660 398414 157140 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 397794 244852 398414 298872 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 397794 368088 398414 410076 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 397794 548640 398414 603728 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 397794 672944 398414 701808 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 433794 2128 434414 157264 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 433794 244852 434414 298996 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 433794 368088 434414 410200 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 433794 548516 434414 603852 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 433794 672944 434414 701808 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 469794 2128 470414 38064 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 469794 122660 470414 157264 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 469794 244852 470414 410200 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 469794 548516 470414 701808 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 505794 2128 506414 37940 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 505794 122660 506414 603728 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 505794 655298 506414 701808 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 541794 2128 542414 38064 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 541794 122660 542414 701808 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 577794 2128 578414 701808 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s 1056 2866 582868 3486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s 1056 38866 582868 39486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s 1056 74866 582868 75486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s 1056 110866 582868 111486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s 1056 146866 582868 147486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s 1056 182866 582868 183486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s 1056 218866 582868 219486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s 1056 254866 582868 255486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s 1056 290866 582868 291486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s 1056 326866 582868 327486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s 1056 362866 582868 363486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s 1056 398866 582868 399486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s 1056 434866 582868 435486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s 1056 470866 582868 471486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s 1056 506866 582868 507486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s 1056 542866 582868 543486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s 1056 578866 582868 579486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s 1056 614866 582868 615486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s 1056 650866 582868 651486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s 1056 686866 582868 687486 6 vccd1
port 532 nsew power bidirectional
rlabel metal5 s 1794 548110 146414 548730 6 vccd1
port 532 nsew power bidirectional
rlabel metal4 s 9234 2128 9854 701808 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 45234 201136 45854 293048 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 81234 201136 81854 293048 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 117234 201260 117854 292924 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 153234 2128 153854 113548 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 153234 201136 153854 293048 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 153234 431364 153854 701808 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 189234 2128 189854 701808 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 225234 2128 225854 701808 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 261234 2128 261854 701808 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 297234 2128 297854 701808 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 333234 122660 333854 701808 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 369234 244976 369854 298872 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 369234 368088 369854 410076 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 369234 548516 369854 603728 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 405234 244852 405854 298872 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 405234 368088 405854 410076 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 405234 548640 405854 603728 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 441234 2128 441854 157264 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 441234 244852 441854 410200 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 441234 548516 441854 701808 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 477234 244852 477854 410200 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 477234 548516 477854 701808 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 513234 122660 513854 701808 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 549234 122660 549854 701808 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s 1056 10306 582868 10926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s 1056 46306 582868 46926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s 1056 82306 582868 82926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s 1056 118306 582868 118926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s 1056 154306 582868 154926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s 1056 190306 582868 190926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s 1056 226306 582868 226926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s 1056 262306 582868 262926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s 1056 298306 582868 298926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s 1056 334306 582868 334926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s 1056 370306 582868 370926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s 1056 406306 582868 406926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s 1056 442306 582868 442926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s 1056 478306 582868 478926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s 1056 514306 582868 514926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s 1056 550306 582868 550926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s 1056 586306 582868 586926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s 1056 622306 582868 622926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s 1056 658306 582868 658926 6 vccd2
port 533 nsew power bidirectional
rlabel metal5 s 1056 694306 582868 694926 6 vccd2
port 533 nsew power bidirectional
rlabel metal4 s 16674 2128 17294 701808 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 52674 201136 53294 293048 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 88674 201136 89294 292924 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 124674 201260 125294 292924 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 160674 2128 161294 113548 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 160674 201260 161294 293048 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 160674 431364 161294 701808 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 196674 2128 197294 701808 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 232674 2128 233294 701808 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 268674 2128 269294 701808 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 304674 2128 305294 701808 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 340674 548516 341294 603852 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 376674 548516 377294 603852 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 412674 548640 413294 603852 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 448674 2128 449294 157264 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 448674 244852 449294 410200 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 448674 548516 449294 701808 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 484674 122784 485294 701808 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 520674 122660 521294 701808 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 556674 2128 557294 701808 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s 1056 17746 582868 18366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s 1056 53746 582868 54366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s 1056 89746 582868 90366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s 1056 125746 582868 126366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s 1056 161746 582868 162366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s 1056 197746 582868 198366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s 1056 233746 582868 234366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s 1056 269746 582868 270366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s 1056 305746 582868 306366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s 1056 341746 582868 342366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s 1056 377746 582868 378366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s 1056 413746 582868 414366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s 1056 449746 582868 450366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s 1056 485746 582868 486366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s 1056 521746 582868 522366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s 1056 557746 582868 558366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s 1056 593746 582868 594366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s 1056 629746 582868 630366 6 vdda1
port 534 nsew power bidirectional
rlabel metal5 s 1056 665746 582868 666366 6 vdda1
port 534 nsew power bidirectional
rlabel metal4 s 24114 2128 24734 701808 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 60114 201136 60734 292924 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 96114 201136 96734 292924 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 132114 201260 132734 292924 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 168114 2128 168734 113548 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 168114 201136 168734 293048 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 168114 431364 168734 701808 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 204114 2128 204734 701808 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 240114 2128 240734 701808 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 276114 2128 276734 701808 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 312114 2128 312734 701808 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 348114 548516 348734 603852 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 384114 548516 384734 603728 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 420114 548640 420734 603852 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 456114 244852 456734 410200 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 456114 548516 456734 701808 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 492114 122660 492734 701808 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 528114 122660 528734 701808 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 564114 2128 564734 701808 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s 1056 25186 582868 25806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s 1056 61186 582868 61806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s 1056 97186 582868 97806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s 1056 133186 582868 133806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s 1056 169186 582868 169806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s 1056 205186 582868 205806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s 1056 241186 582868 241806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s 1056 277186 582868 277806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s 1056 313186 582868 313806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s 1056 349186 582868 349806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s 1056 385186 582868 385806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s 1056 421186 582868 421806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s 1056 457186 582868 457806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s 1056 493186 582868 493806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s 1056 529186 582868 529806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s 1056 565186 582868 565806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s 1056 601186 582868 601806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s 1056 637186 582868 637806 6 vdda2
port 535 nsew power bidirectional
rlabel metal5 s 1056 673186 582868 673806 6 vdda2
port 535 nsew power bidirectional
rlabel metal4 s 20394 2128 21014 701808 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 56394 201136 57014 292924 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 92394 201260 93014 292924 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 128394 201136 129014 293048 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 164394 2128 165014 113548 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 164394 201136 165014 293048 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 164394 431364 165014 701808 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 200394 2128 201014 701808 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 236394 2128 237014 701808 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 272394 2128 273014 701808 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 308394 2128 309014 701808 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 344394 548516 345014 603852 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 380394 548640 381014 603728 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 416394 548516 417014 603852 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 452394 2128 453014 157264 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 452394 244852 453014 410200 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 452394 548516 453014 701808 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 488394 122660 489014 701808 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 524394 122660 525014 701808 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 560394 2128 561014 701808 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s 1056 21466 582868 22086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s 1056 57466 582868 58086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s 1056 93466 582868 94086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s 1056 129466 582868 130086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s 1056 165466 582868 166086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s 1056 201466 582868 202086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s 1056 237466 582868 238086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s 1056 273466 582868 274086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s 1056 309466 582868 310086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s 1056 345466 582868 346086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s 1056 381466 582868 382086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s 1056 417466 582868 418086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s 1056 453466 582868 454086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s 1056 489466 582868 490086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s 1056 525466 582868 526086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s 1056 561466 582868 562086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s 1056 597466 582868 598086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s 1056 633466 582868 634086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal5 s 1056 669466 582868 670086 6 vssa1
port 536 nsew ground bidirectional
rlabel metal4 s 27834 2128 28454 701808 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 63834 201136 64454 292924 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 99834 201260 100454 292924 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 135834 201136 136454 293048 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 135834 546808 136454 701808 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 171834 2128 172454 113548 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 171834 201136 172454 293048 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 171834 431364 172454 701808 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 207834 2128 208454 701808 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 243834 2128 244454 701808 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 279834 2128 280454 701808 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 315834 2128 316454 701808 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 351834 244852 352454 298996 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 387834 244852 388454 298872 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 423834 2128 424454 157264 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 423834 244852 424454 298872 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 459834 244852 460454 410200 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 459834 548516 460454 701808 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 495834 122660 496454 701808 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 531834 122660 532454 701808 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 567834 2128 568454 701808 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s 1056 28906 582868 29526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s 1056 64906 582868 65526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s 1056 100906 582868 101526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s 1056 136906 582868 137526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s 1056 172906 582868 173526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s 1056 208906 582868 209526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s 1056 244906 582868 245526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s 1056 280906 582868 281526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s 1056 316906 582868 317526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s 1056 352906 582868 353526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s 1056 388906 582868 389526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s 1056 424906 582868 425526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s 1056 460906 582868 461526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s 1056 496906 582868 497526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s 1056 532906 582868 533526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s 1056 568906 582868 569526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s 1056 604906 582868 605526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s 1056 640906 582868 641526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal5 s 1056 676906 582868 677526 6 vssa2
port 537 nsew ground bidirectional
rlabel metal4 s 5514 2128 6134 701808 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 41514 2128 42134 33464 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 41514 82020 42134 113548 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 41514 201136 42134 293048 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 41514 431364 42134 462212 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 41514 546808 42134 577112 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 41514 670412 42134 701808 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 77514 2128 78134 33340 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 77514 82020 78134 113424 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 77514 201260 78134 292924 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 77514 431488 78134 462088 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 77514 546808 78134 577112 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 77514 670412 78134 701808 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 113514 2128 114134 33464 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 113514 82020 114134 113548 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 113514 201136 114134 293048 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 113514 431364 114134 462212 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 113514 546808 114134 577112 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 113514 670412 114134 701808 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 149514 2128 150134 113548 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 149514 201136 150134 293048 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 149514 431364 150134 701808 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 185514 2128 186134 701808 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 221514 2128 222134 701808 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 257514 2128 258134 701808 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 293514 2128 294134 701808 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 329514 2128 330134 38064 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 329514 122660 330134 701808 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 365514 2128 366134 37940 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 365514 122784 366134 157140 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 365514 244852 366134 298872 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 365514 368088 366134 410076 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 365514 548516 366134 603728 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 365514 672944 366134 701808 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 401514 2128 402134 38064 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 401514 122784 402134 157264 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 401514 244852 402134 298872 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 401514 368088 402134 410200 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 401514 548516 402134 603728 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 401514 672944 402134 701808 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 437514 2128 438134 157264 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 437514 244852 438134 298996 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 437514 368088 438134 410076 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 437514 548640 438134 603852 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 437514 672944 438134 701808 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 473514 2128 474134 37940 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 473514 122660 474134 157264 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 473514 244852 474134 410200 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 473514 548640 474134 701808 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 509514 2128 510134 38064 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 509514 122660 510134 701808 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 545514 2128 546134 38064 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 545514 122660 546134 701808 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 581514 2128 582134 701808 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s 1056 6586 582868 7206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s 1056 42586 582868 43206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s 1056 78586 582868 79206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s 1056 114586 582868 115206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s 1056 150586 582868 151206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s 1056 186586 582868 187206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s 1056 222586 582868 223206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s 1056 258586 582868 259206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s 1056 294586 582868 295206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s 1056 330586 582868 331206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s 1056 366586 582868 367206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s 1056 402586 582868 403206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s 1056 438586 582868 439206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s 1056 474586 582868 475206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s 1056 510586 582868 511206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s 1056 546586 582868 547206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s 1056 582586 582868 583206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s 1056 618586 582868 619206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s 1056 654586 582868 655206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s 1056 690586 582868 691206 6 vssd1
port 538 nsew ground bidirectional
rlabel metal5 s 5514 83670 150134 84290 6 vssd1
port 538 nsew ground bidirectional
rlabel metal4 s 12954 2128 13574 701808 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 48954 201136 49574 293048 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 84954 201260 85574 292924 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 120954 201136 121574 293048 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 156954 2128 157574 113548 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 156954 201136 157574 293048 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 156954 431364 157574 701808 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 192954 2128 193574 701808 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 228954 2128 229574 701808 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 264954 2128 265574 701808 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 300954 2128 301574 701808 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 336954 122660 337574 701808 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 372954 368088 373574 410076 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 372954 548640 373574 603852 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 408954 368088 409574 410200 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 408954 548516 409574 603852 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 444954 2128 445574 157264 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 444954 244852 445574 410076 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 444954 548640 445574 701808 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 480954 122660 481574 410200 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 480954 548516 481574 701808 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 516954 122660 517574 701808 6 vssd2
port 539 nsew ground bidirectional
rlabel metal4 s 552954 122660 553574 701808 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s 1056 14026 582868 14646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s 1056 50026 582868 50646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s 1056 86026 582868 86646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s 1056 122026 582868 122646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s 1056 158026 582868 158646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s 1056 194026 582868 194646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s 1056 230026 582868 230646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s 1056 266026 582868 266646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s 1056 302026 582868 302646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s 1056 338026 582868 338646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s 1056 374026 582868 374646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s 1056 410026 582868 410646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s 1056 446026 582868 446646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s 1056 482026 582868 482646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s 1056 518026 582868 518646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s 1056 554026 582868 554646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s 1056 590026 582868 590646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s 1056 626026 582868 626646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s 1056 662026 582868 662646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal5 s 1056 698026 582868 698646 6 vssd2
port 539 nsew ground bidirectional
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 540 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 541 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 542 nsew signal output
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 543 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 544 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 545 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 546 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 547 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 548 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 549 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 550 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 551 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 552 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 553 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 554 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 555 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 556 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 557 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 558 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 559 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 560 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 561 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 562 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 563 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 564 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 565 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 566 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 567 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 568 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 569 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 570 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 571 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 572 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 573 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 574 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 575 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 576 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 577 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 578 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 579 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 580 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 581 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 582 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 583 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 584 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 585 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 586 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 587 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 588 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 589 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 590 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 591 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 592 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 593 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 594 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 595 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 596 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 597 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 598 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 599 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 600 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 601 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 602 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 603 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 604 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 605 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 606 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 607 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 608 nsew signal output
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 609 nsew signal output
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 610 nsew signal output
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 611 nsew signal output
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 612 nsew signal output
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 613 nsew signal output
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 614 nsew signal output
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 615 nsew signal output
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 616 nsew signal output
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 617 nsew signal output
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 618 nsew signal output
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 619 nsew signal output
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 620 nsew signal output
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 621 nsew signal output
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 622 nsew signal output
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 623 nsew signal output
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 624 nsew signal output
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 625 nsew signal output
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 626 nsew signal output
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 627 nsew signal output
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 628 nsew signal output
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 629 nsew signal output
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 630 nsew signal output
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 631 nsew signal output
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 632 nsew signal output
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 633 nsew signal output
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 634 nsew signal output
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 635 nsew signal output
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 636 nsew signal output
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 637 nsew signal output
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 638 nsew signal output
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 639 nsew signal output
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 640 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 641 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 642 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 643 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 644 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 645 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 174174288
string GDS_FILE /home/mkhan33/mpw8/openram_testchip2/openlane/user_project_wrapper/runs/22_12_19_00_13/results/signoff/user_project_wrapper.magic.gds
string GDS_START 70228282
<< end >>


VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO rram_test
  CLASS BLOCK ;
  FOREIGN rram_test ;
  ORIGIN 12.990 16.000 ;
  SIZE 42.870 BY 23.350 ;
  PIN RE_BR0
    ANTENNADIFFAREA 4.200000 ;
    PORT
      LAYER li1 ;
        RECT 12.075 -2.820 12.245 2.530 ;
        RECT 12.075 -12.820 12.245 -7.470 ;
      LAYER mcon ;
        RECT 12.075 2.145 12.245 2.315 ;
        RECT 12.075 1.785 12.245 1.955 ;
        RECT 12.075 1.425 12.245 1.595 ;
        RECT 12.075 1.065 12.245 1.235 ;
        RECT 12.075 0.705 12.245 0.875 ;
        RECT 12.075 0.345 12.245 0.515 ;
        RECT 12.075 -0.015 12.245 0.155 ;
        RECT 12.075 -0.375 12.245 -0.205 ;
        RECT 12.075 -0.735 12.245 -0.565 ;
        RECT 12.075 -1.095 12.245 -0.925 ;
        RECT 12.075 -1.455 12.245 -1.285 ;
        RECT 12.075 -1.815 12.245 -1.645 ;
        RECT 12.075 -2.175 12.245 -2.005 ;
        RECT 12.075 -2.535 12.245 -2.365 ;
        RECT 12.075 -7.855 12.245 -7.685 ;
        RECT 12.075 -8.215 12.245 -8.045 ;
        RECT 12.075 -8.575 12.245 -8.405 ;
        RECT 12.075 -8.935 12.245 -8.765 ;
        RECT 12.075 -9.295 12.245 -9.125 ;
        RECT 12.075 -9.655 12.245 -9.485 ;
        RECT 12.075 -10.015 12.245 -9.845 ;
        RECT 12.075 -10.375 12.245 -10.205 ;
        RECT 12.075 -10.735 12.245 -10.565 ;
        RECT 12.075 -11.095 12.245 -10.925 ;
        RECT 12.075 -11.455 12.245 -11.285 ;
        RECT 12.075 -11.815 12.245 -11.645 ;
        RECT 12.075 -12.175 12.245 -12.005 ;
        RECT 12.075 -12.535 12.245 -12.365 ;
      LAYER met1 ;
        RECT 12.030 -3.080 12.350 2.535 ;
        RECT 12.030 -3.285 14.945 -3.080 ;
        RECT 14.665 -4.970 14.945 -3.285 ;
        RECT 12.030 -13.080 12.350 -7.465 ;
        RECT 12.030 -13.285 14.945 -13.080 ;
        RECT 14.665 -14.970 14.945 -13.285 ;
      LAYER via ;
        RECT 12.060 2.070 12.320 2.330 ;
        RECT 12.060 1.750 12.320 2.010 ;
        RECT 12.060 1.430 12.320 1.690 ;
        RECT 12.060 1.110 12.320 1.370 ;
        RECT 12.060 0.790 12.320 1.050 ;
        RECT 12.060 0.470 12.320 0.730 ;
        RECT 12.060 0.150 12.320 0.410 ;
        RECT 12.060 -0.170 12.320 0.090 ;
        RECT 12.060 -0.490 12.320 -0.230 ;
        RECT 12.060 -0.810 12.320 -0.550 ;
        RECT 12.060 -1.130 12.320 -0.870 ;
        RECT 12.060 -1.450 12.320 -1.190 ;
        RECT 12.060 -1.770 12.320 -1.510 ;
        RECT 12.060 -2.090 12.320 -1.830 ;
        RECT 12.060 -2.410 12.320 -2.150 ;
        RECT 12.060 -2.730 12.320 -2.470 ;
        RECT 14.670 -4.910 14.930 -4.650 ;
        RECT 12.060 -7.930 12.320 -7.670 ;
        RECT 12.060 -8.250 12.320 -7.990 ;
        RECT 12.060 -8.570 12.320 -8.310 ;
        RECT 12.060 -8.890 12.320 -8.630 ;
        RECT 12.060 -9.210 12.320 -8.950 ;
        RECT 12.060 -9.530 12.320 -9.270 ;
        RECT 12.060 -9.850 12.320 -9.590 ;
        RECT 12.060 -10.170 12.320 -9.910 ;
        RECT 12.060 -10.490 12.320 -10.230 ;
        RECT 12.060 -10.810 12.320 -10.550 ;
        RECT 12.060 -11.130 12.320 -10.870 ;
        RECT 12.060 -11.450 12.320 -11.190 ;
        RECT 12.060 -11.770 12.320 -11.510 ;
        RECT 12.060 -12.090 12.320 -11.830 ;
        RECT 12.060 -12.410 12.320 -12.150 ;
        RECT 12.060 -12.730 12.320 -12.470 ;
        RECT 14.670 -14.910 14.930 -14.650 ;
      LAYER met2 ;
        RECT 12.425 5.570 14.240 7.350 ;
        RECT 13.910 5.220 14.240 5.570 ;
        RECT 13.910 4.990 14.950 5.220 ;
        RECT 12.030 -2.815 12.350 2.535 ;
        RECT 14.445 -4.580 14.950 4.990 ;
        RECT 12.030 -12.815 12.350 -7.465 ;
        RECT 14.440 -14.970 14.945 -4.580 ;
        RECT 14.435 -16.000 14.940 -14.970 ;
    END
  END RE_BR0
  PIN WL0
    ANTENNAGATEAREA 0.216000 ;
    PORT
      LAYER li1 ;
        RECT 8.640 -3.615 8.955 -3.060 ;
        RECT 18.640 -3.615 18.955 -3.060 ;
        RECT 25.270 -3.615 25.670 -3.365 ;
        RECT 7.635 -3.785 25.670 -3.615 ;
      LAYER mcon ;
        RECT 25.375 -3.660 25.545 -3.490 ;
      LAYER met1 ;
        RECT 25.270 -3.785 25.670 -3.365 ;
      LAYER via ;
        RECT 25.345 -3.700 25.605 -3.440 ;
      LAYER met2 ;
        RECT 22.200 5.570 24.015 7.350 ;
        RECT 23.605 4.695 24.010 5.570 ;
        RECT 23.605 4.535 25.670 4.695 ;
        RECT 25.270 -3.785 25.670 4.535 ;
    END
  END WL0
  PIN WL1
    ANTENNAGATEAREA 0.216000 ;
    PORT
      LAYER li1 ;
        RECT 8.640 -13.615 8.955 -13.060 ;
        RECT 18.640 -13.615 18.955 -13.060 ;
        RECT 26.820 -13.615 27.220 -13.325 ;
        RECT 7.635 -13.785 27.220 -13.615 ;
      LAYER mcon ;
        RECT 26.925 -13.620 27.095 -13.450 ;
      LAYER met1 ;
        RECT 26.820 -13.745 27.220 -13.325 ;
      LAYER via ;
        RECT 26.895 -13.660 27.155 -13.400 ;
      LAYER met2 ;
        RECT 26.110 5.570 27.925 7.350 ;
        RECT 26.820 -13.745 27.220 5.570 ;
    END
  END WL1
  PIN RE_WL0
    ANTENNAGATEAREA 4.200000 ;
    PORT
      LAYER li1 ;
        RECT 25.970 -4.075 26.370 -3.825 ;
        RECT 7.635 -4.245 26.370 -4.075 ;
        RECT 7.980 -4.925 8.335 -4.245 ;
        RECT 12.255 -4.925 12.610 -4.245 ;
        RECT 17.980 -4.925 18.335 -4.245 ;
        RECT 22.255 -4.925 22.610 -4.245 ;
      LAYER mcon ;
        RECT 26.075 -4.120 26.245 -3.950 ;
      LAYER met1 ;
        RECT 25.970 -4.245 26.370 -3.825 ;
      LAYER via ;
        RECT 26.045 -4.160 26.305 -3.900 ;
      LAYER met2 ;
        RECT 24.155 5.570 25.970 7.350 ;
        RECT 25.590 5.270 25.970 5.570 ;
        RECT 25.590 4.910 26.370 5.270 ;
        RECT 25.970 -4.245 26.370 4.910 ;
    END
  END RE_WL0
  PIN RE_WL1
    ANTENNAGATEAREA 4.200000 ;
    PORT
      LAYER li1 ;
        RECT 28.380 -14.075 28.780 -13.825 ;
        RECT 7.635 -14.245 28.780 -14.075 ;
        RECT 7.980 -14.925 8.335 -14.245 ;
        RECT 12.255 -14.925 12.610 -14.245 ;
        RECT 17.980 -14.925 18.335 -14.245 ;
        RECT 22.255 -14.925 22.610 -14.245 ;
      LAYER mcon ;
        RECT 28.485 -14.120 28.655 -13.950 ;
      LAYER met1 ;
        RECT 28.380 -14.245 28.780 -13.825 ;
      LAYER via ;
        RECT 28.455 -14.160 28.715 -13.900 ;
      LAYER met2 ;
        RECT 28.065 5.570 29.880 7.350 ;
        RECT 28.380 -14.245 28.780 5.570 ;
    END
  END RE_WL1
  PIN VDD
    ANTENNADIFFAREA 0.905600 ;
    PORT
      LAYER li1 ;
        RECT 9.145 -0.590 9.395 -0.260 ;
        RECT 19.145 -0.590 19.395 -0.260 ;
        RECT 9.165 -2.505 9.425 -1.925 ;
        RECT 19.165 -2.505 19.425 -1.925 ;
        RECT 9.145 -10.590 9.395 -10.260 ;
        RECT 19.145 -10.590 19.395 -10.260 ;
        RECT 9.165 -12.505 9.425 -11.925 ;
        RECT 19.165 -12.505 19.425 -11.925 ;
      LAYER mcon ;
        RECT 9.225 -0.510 9.395 -0.340 ;
        RECT 19.225 -0.510 19.395 -0.340 ;
        RECT 9.215 -2.360 9.385 -2.190 ;
        RECT 19.215 -2.360 19.385 -2.190 ;
        RECT 9.225 -10.510 9.395 -10.340 ;
        RECT 19.225 -10.510 19.395 -10.340 ;
        RECT 9.215 -12.360 9.385 -12.190 ;
        RECT 19.215 -12.360 19.385 -12.190 ;
      LAYER met1 ;
        RECT 5.485 4.875 18.110 5.220 ;
        RECT 9.165 0.360 9.425 0.780 ;
        RECT 19.165 0.360 19.425 0.780 ;
        RECT 9.165 0.040 9.485 0.360 ;
        RECT 19.165 0.040 19.485 0.360 ;
        RECT 9.165 -0.280 9.425 0.040 ;
        RECT 19.165 -0.280 19.425 0.040 ;
        RECT 9.165 -0.570 9.455 -0.280 ;
        RECT 19.165 -0.570 19.455 -0.280 ;
        RECT 6.690 -3.855 7.050 -3.685 ;
        RECT 9.165 -3.855 9.425 -0.570 ;
        RECT 6.690 -4.060 9.425 -3.855 ;
        RECT 16.690 -3.855 17.050 -3.685 ;
        RECT 19.165 -3.855 19.425 -0.570 ;
        RECT 16.690 -4.060 19.425 -3.855 ;
        RECT 9.165 -9.640 9.425 -9.220 ;
        RECT 19.165 -9.640 19.425 -9.220 ;
        RECT 9.165 -9.960 9.485 -9.640 ;
        RECT 19.165 -9.960 19.485 -9.640 ;
        RECT 9.165 -10.280 9.425 -9.960 ;
        RECT 19.165 -10.280 19.425 -9.960 ;
        RECT 9.165 -10.570 9.455 -10.280 ;
        RECT 19.165 -10.570 19.455 -10.280 ;
        RECT 6.690 -13.855 7.050 -13.685 ;
        RECT 9.165 -13.855 9.425 -10.570 ;
        RECT 6.690 -14.060 9.425 -13.855 ;
        RECT 16.690 -13.855 17.050 -13.685 ;
        RECT 19.165 -13.855 19.425 -10.570 ;
        RECT 16.690 -14.060 19.425 -13.855 ;
      LAYER via ;
        RECT 6.730 4.910 6.990 5.170 ;
        RECT 17.495 4.910 17.755 5.170 ;
        RECT 9.195 0.070 9.455 0.330 ;
        RECT 19.195 0.070 19.455 0.330 ;
        RECT 6.735 -3.995 6.995 -3.735 ;
        RECT 16.735 -3.995 16.995 -3.735 ;
        RECT 9.195 -9.930 9.455 -9.670 ;
        RECT 19.195 -9.930 19.455 -9.670 ;
        RECT 6.735 -13.995 6.995 -13.735 ;
        RECT 16.735 -13.995 16.995 -13.735 ;
      LAYER met2 ;
        RECT 6.560 5.570 8.375 7.350 ;
        RECT 6.690 -16.000 7.055 5.570 ;
        RECT 17.055 4.760 18.110 5.320 ;
        RECT 16.685 4.450 18.110 4.760 ;
        RECT 9.145 0.040 11.015 0.360 ;
        RECT 16.685 -3.680 17.055 4.450 ;
        RECT 19.145 0.040 21.015 0.360 ;
        RECT 9.145 -9.960 11.015 -9.640 ;
        RECT 16.690 -16.000 17.055 -3.680 ;
        RECT 19.145 -9.960 21.015 -9.640 ;
    END
  END VDD
  PIN p036_SL
    ANTENNAGATEAREA 0.054000 ;
    PORT
      LAYER li1 ;
        RECT 0.730 1.505 1.290 1.790 ;
      LAYER mcon ;
        RECT 1.065 1.555 1.235 1.725 ;
      LAYER met1 ;
        RECT 0.930 1.505 1.365 1.790 ;
      LAYER via ;
        RECT 1.015 1.530 1.275 1.790 ;
      LAYER met2 ;
        RECT -7.125 5.570 -5.310 7.350 ;
        RECT -5.760 1.790 -5.455 5.570 ;
        RECT -5.760 1.515 1.370 1.790 ;
    END
  END p036_SL
  PIN p700_SL
    ANTENNAGATEAREA 1.050000 ;
    PORT
      LAYER li1 ;
        RECT 4.045 -5.105 4.400 -4.820 ;
      LAYER mcon ;
        RECT 4.135 -5.025 4.305 -4.855 ;
      LAYER met1 ;
        RECT 3.890 -5.225 4.555 -4.655 ;
      LAYER via ;
        RECT 4.085 -5.065 4.345 -4.805 ;
      LAYER met2 ;
        RECT -12.990 5.570 -11.175 7.350 ;
        RECT -11.795 -4.810 -11.320 5.570 ;
        RECT 3.900 -4.810 4.560 -4.655 ;
        RECT -11.795 -5.100 4.710 -4.810 ;
        RECT 3.900 -5.230 4.560 -5.100 ;
    END
  END p700_SL
  PIN p300_SL
    ANTENNAGATEAREA 0.450000 ;
    PORT
      LAYER li1 ;
        RECT 2.995 -1.095 3.555 -0.810 ;
      LAYER mcon ;
        RECT 3.330 -1.045 3.500 -0.875 ;
      LAYER met1 ;
        RECT 3.195 -1.095 3.630 -0.810 ;
      LAYER via ;
        RECT 3.280 -1.070 3.540 -0.810 ;
      LAYER met2 ;
        RECT -11.035 5.570 -9.220 7.350 ;
        RECT -9.840 -0.815 -9.365 5.570 ;
        RECT 3.195 -0.815 3.630 -0.810 ;
        RECT -9.840 -1.085 3.630 -0.815 ;
    END
  END p300_SL
  PIN p100_SL
    ANTENNAGATEAREA 0.150000 ;
    PORT
      LAYER li1 ;
        RECT 1.945 0.740 2.505 1.025 ;
      LAYER mcon ;
        RECT 2.280 0.790 2.450 0.960 ;
      LAYER met1 ;
        RECT 2.145 0.740 2.580 1.025 ;
      LAYER via ;
        RECT 2.230 0.765 2.490 1.025 ;
      LAYER met2 ;
        RECT -9.080 5.570 -7.265 7.350 ;
        RECT -7.885 1.030 -7.510 5.570 ;
        RECT -7.885 0.755 2.590 1.030 ;
    END
  END p100_SL
  PIN p1T1R_WL
    ANTENNADIFFAREA 3.408000 ;
    PORT
      LAYER li1 ;
        RECT 0.560 2.020 0.730 2.350 ;
        RECT 1.775 1.400 1.945 2.350 ;
        RECT 2.830 -0.635 3.000 2.350 ;
        RECT 3.865 -3.000 4.035 2.350 ;
      LAYER mcon ;
        RECT 0.560 2.100 0.730 2.270 ;
        RECT 1.775 1.980 1.945 2.150 ;
        RECT 1.775 1.620 1.945 1.790 ;
        RECT 2.830 1.800 3.000 1.970 ;
        RECT 2.830 1.440 3.000 1.610 ;
        RECT 2.830 1.080 3.000 1.250 ;
        RECT 2.830 0.720 3.000 0.890 ;
        RECT 2.830 0.360 3.000 0.530 ;
        RECT 2.830 0.000 3.000 0.170 ;
        RECT 2.830 -0.360 3.000 -0.190 ;
        RECT 3.865 1.965 4.035 2.135 ;
        RECT 3.865 1.605 4.035 1.775 ;
        RECT 3.865 1.245 4.035 1.415 ;
        RECT 3.865 0.885 4.035 1.055 ;
        RECT 3.865 0.525 4.035 0.695 ;
        RECT 3.865 0.165 4.035 0.335 ;
        RECT 3.865 -0.195 4.035 -0.025 ;
        RECT 3.865 -0.555 4.035 -0.385 ;
        RECT 3.865 -0.915 4.035 -0.745 ;
        RECT 3.865 -1.275 4.035 -1.105 ;
        RECT 3.865 -1.635 4.035 -1.465 ;
        RECT 3.865 -1.995 4.035 -1.825 ;
        RECT 3.865 -2.355 4.035 -2.185 ;
        RECT 3.865 -2.715 4.035 -2.545 ;
      LAYER met1 ;
        RECT 0.515 2.035 0.835 2.355 ;
        RECT 1.730 1.395 2.050 2.355 ;
        RECT 2.785 -0.635 3.105 2.355 ;
        RECT 3.820 -3.000 4.140 2.355 ;
      LAYER via ;
        RECT 0.545 2.065 0.805 2.325 ;
        RECT 1.760 1.915 2.020 2.175 ;
        RECT 1.760 1.595 2.020 1.855 ;
        RECT 2.815 1.810 3.075 2.070 ;
        RECT 2.815 1.490 3.075 1.750 ;
        RECT 2.815 1.170 3.075 1.430 ;
        RECT 2.815 0.850 3.075 1.110 ;
        RECT 2.815 0.530 3.075 0.790 ;
        RECT 2.815 0.210 3.075 0.470 ;
        RECT 2.815 -0.110 3.075 0.150 ;
        RECT 2.815 -0.430 3.075 -0.170 ;
        RECT 3.850 1.890 4.110 2.150 ;
        RECT 3.850 1.570 4.110 1.830 ;
        RECT 3.850 1.250 4.110 1.510 ;
        RECT 3.850 0.930 4.110 1.190 ;
        RECT 3.850 0.610 4.110 0.870 ;
        RECT 3.850 0.290 4.110 0.550 ;
        RECT 3.850 -0.030 4.110 0.230 ;
        RECT 3.850 -0.350 4.110 -0.090 ;
        RECT 3.850 -0.670 4.110 -0.410 ;
        RECT 3.850 -0.990 4.110 -0.730 ;
        RECT 3.850 -1.310 4.110 -1.050 ;
        RECT 3.850 -1.630 4.110 -1.370 ;
        RECT 3.850 -1.950 4.110 -1.690 ;
        RECT 3.850 -2.270 4.110 -2.010 ;
        RECT 3.850 -2.590 4.110 -2.330 ;
        RECT 3.850 -2.910 4.110 -2.650 ;
      LAYER met2 ;
        RECT -5.170 5.570 -3.355 7.350 ;
        RECT -3.860 2.355 -3.560 5.570 ;
        RECT -3.860 2.035 4.140 2.355 ;
        RECT 1.730 1.395 2.050 2.035 ;
        RECT 2.785 -0.565 3.105 2.035 ;
        RECT 3.820 -2.995 4.140 2.035 ;
    END
  END p1T1R_WL
  PIN p1T1R_TE
    ANTENNADIFFAREA 3.408000 ;
    PORT
      LAYER li1 ;
        RECT 1.060 2.020 1.230 2.350 ;
        RECT 2.275 1.400 2.445 2.350 ;
        RECT 3.330 -0.635 3.500 2.350 ;
        RECT 4.365 -3.000 4.535 2.350 ;
      LAYER mcon ;
        RECT 1.060 2.100 1.230 2.270 ;
        RECT 2.275 1.975 2.445 2.145 ;
        RECT 2.275 1.615 2.445 1.785 ;
        RECT 3.330 1.800 3.500 1.970 ;
        RECT 3.330 1.440 3.500 1.610 ;
        RECT 3.330 1.080 3.500 1.250 ;
        RECT 3.330 0.720 3.500 0.890 ;
        RECT 3.330 0.360 3.500 0.530 ;
        RECT 3.330 0.000 3.500 0.170 ;
        RECT 3.330 -0.360 3.500 -0.190 ;
        RECT 4.365 1.960 4.535 2.130 ;
        RECT 4.365 1.600 4.535 1.770 ;
        RECT 4.365 1.240 4.535 1.410 ;
        RECT 4.365 0.880 4.535 1.050 ;
        RECT 4.365 0.520 4.535 0.690 ;
        RECT 4.365 0.160 4.535 0.330 ;
        RECT 4.365 -0.200 4.535 -0.030 ;
        RECT 4.365 -0.560 4.535 -0.390 ;
        RECT 4.365 -0.920 4.535 -0.750 ;
        RECT 4.365 -1.280 4.535 -1.110 ;
        RECT 4.365 -1.640 4.535 -1.470 ;
        RECT 4.365 -2.000 4.535 -1.830 ;
        RECT 4.365 -2.360 4.535 -2.190 ;
        RECT 4.365 -2.720 4.535 -2.550 ;
      LAYER met1 ;
        RECT 0.720 2.950 1.040 3.210 ;
        RECT 1.935 2.950 2.255 3.210 ;
        RECT 2.990 2.950 3.310 3.210 ;
        RECT 4.025 2.950 4.345 3.210 ;
        RECT 0.820 2.635 0.980 2.950 ;
        RECT 2.035 2.635 2.195 2.950 ;
        RECT 3.090 2.635 3.250 2.950 ;
        RECT 4.125 2.635 4.285 2.950 ;
        RECT 0.820 2.495 1.215 2.635 ;
        RECT 2.035 2.495 2.430 2.635 ;
        RECT 3.090 2.495 3.485 2.635 ;
        RECT 4.125 2.495 4.520 2.635 ;
        RECT 1.075 2.330 1.215 2.495 ;
        RECT 2.290 2.330 2.430 2.495 ;
        RECT 3.345 2.330 3.485 2.495 ;
        RECT 4.380 2.330 4.520 2.495 ;
        RECT 1.030 2.020 1.260 2.330 ;
        RECT 2.245 1.395 2.475 2.330 ;
        RECT 3.300 -0.635 3.530 2.330 ;
        RECT 4.335 -3.000 4.565 2.330 ;
      LAYER via ;
        RECT 0.750 2.950 1.010 3.210 ;
        RECT 1.965 2.950 2.225 3.210 ;
        RECT 3.020 2.950 3.280 3.210 ;
        RECT 4.055 2.950 4.315 3.210 ;
      LAYER met2 ;
        RECT -3.215 5.570 -1.400 7.350 ;
        RECT -1.815 3.245 -1.400 5.570 ;
        RECT -1.815 2.900 4.390 3.245 ;
    END
  END p1T1R_TE
  PIN p1R_SL
    PORT
      LAYER met1 ;
        RECT -0.460 4.435 0.840 4.695 ;
      LAYER via ;
        RECT -0.420 4.435 -0.160 4.695 ;
        RECT 0.550 4.435 0.810 4.695 ;
      LAYER met2 ;
        RECT -1.260 5.570 0.555 7.350 ;
        RECT 0.695 5.570 2.510 7.350 ;
        RECT -0.750 4.300 0.195 5.570 ;
        RECT 0.695 4.725 1.250 5.570 ;
        RECT 0.550 4.405 1.250 4.725 ;
    END
  END p1R_SL
  PIN RE_BL0
    ANTENNADIFFAREA 4.200000 ;
    PORT
      LAYER li1 ;
        RECT 7.800 -2.820 7.970 2.530 ;
        RECT 7.800 -12.820 7.970 -7.470 ;
      LAYER mcon ;
        RECT 7.800 2.145 7.970 2.315 ;
        RECT 7.800 1.785 7.970 1.955 ;
        RECT 7.800 1.425 7.970 1.595 ;
        RECT 7.800 1.065 7.970 1.235 ;
        RECT 7.800 0.705 7.970 0.875 ;
        RECT 7.800 0.345 7.970 0.515 ;
        RECT 7.800 -0.015 7.970 0.155 ;
        RECT 7.800 -0.375 7.970 -0.205 ;
        RECT 7.800 -0.735 7.970 -0.565 ;
        RECT 7.800 -1.095 7.970 -0.925 ;
        RECT 7.800 -1.455 7.970 -1.285 ;
        RECT 7.800 -1.815 7.970 -1.645 ;
        RECT 7.800 -2.175 7.970 -2.005 ;
        RECT 7.800 -2.535 7.970 -2.365 ;
        RECT 7.800 -7.855 7.970 -7.685 ;
        RECT 7.800 -8.215 7.970 -8.045 ;
        RECT 7.800 -8.575 7.970 -8.405 ;
        RECT 7.800 -8.935 7.970 -8.765 ;
        RECT 7.800 -9.295 7.970 -9.125 ;
        RECT 7.800 -9.655 7.970 -9.485 ;
        RECT 7.800 -10.015 7.970 -9.845 ;
        RECT 7.800 -10.375 7.970 -10.205 ;
        RECT 7.800 -10.735 7.970 -10.565 ;
        RECT 7.800 -11.095 7.970 -10.925 ;
        RECT 7.800 -11.455 7.970 -11.285 ;
        RECT 7.800 -11.815 7.970 -11.645 ;
        RECT 7.800 -12.175 7.970 -12.005 ;
        RECT 7.800 -12.535 7.970 -12.365 ;
      LAYER met1 ;
        RECT 7.755 -2.465 8.075 2.535 ;
        RECT 5.495 -2.780 8.075 -2.465 ;
        RECT 5.495 -4.925 5.860 -2.780 ;
        RECT 7.755 -2.820 8.075 -2.780 ;
        RECT 7.755 -12.465 8.075 -7.465 ;
        RECT 5.495 -12.780 8.075 -12.465 ;
        RECT 5.495 -14.925 5.860 -12.780 ;
        RECT 7.755 -12.820 8.075 -12.780 ;
      LAYER via ;
        RECT 7.785 2.070 8.045 2.330 ;
        RECT 7.785 1.750 8.045 2.010 ;
        RECT 7.785 1.430 8.045 1.690 ;
        RECT 7.785 1.110 8.045 1.370 ;
        RECT 7.785 0.790 8.045 1.050 ;
        RECT 7.785 0.470 8.045 0.730 ;
        RECT 7.785 0.150 8.045 0.410 ;
        RECT 7.785 -0.170 8.045 0.090 ;
        RECT 7.785 -0.490 8.045 -0.230 ;
        RECT 7.785 -0.810 8.045 -0.550 ;
        RECT 7.785 -1.130 8.045 -0.870 ;
        RECT 7.785 -1.450 8.045 -1.190 ;
        RECT 7.785 -1.770 8.045 -1.510 ;
        RECT 7.785 -2.090 8.045 -1.830 ;
        RECT 7.785 -2.410 8.045 -2.150 ;
        RECT 7.785 -2.730 8.045 -2.470 ;
        RECT 5.565 -4.910 5.825 -4.650 ;
        RECT 7.785 -7.930 8.045 -7.670 ;
        RECT 7.785 -8.250 8.045 -7.990 ;
        RECT 7.785 -8.570 8.045 -8.310 ;
        RECT 7.785 -8.890 8.045 -8.630 ;
        RECT 7.785 -9.210 8.045 -8.950 ;
        RECT 7.785 -9.530 8.045 -9.270 ;
        RECT 7.785 -9.850 8.045 -9.590 ;
        RECT 7.785 -10.170 8.045 -9.910 ;
        RECT 7.785 -10.490 8.045 -10.230 ;
        RECT 7.785 -10.810 8.045 -10.550 ;
        RECT 7.785 -11.130 8.045 -10.870 ;
        RECT 7.785 -11.450 8.045 -11.190 ;
        RECT 7.785 -11.770 8.045 -11.510 ;
        RECT 7.785 -12.090 8.045 -11.830 ;
        RECT 7.785 -12.410 8.045 -12.150 ;
        RECT 7.785 -12.730 8.045 -12.470 ;
        RECT 5.565 -14.910 5.825 -14.650 ;
      LAYER met2 ;
        RECT 2.650 5.570 4.465 7.350 ;
        RECT 4.150 5.220 4.465 5.570 ;
        RECT 4.150 4.865 5.990 5.220 ;
        RECT 5.485 -16.000 5.990 4.865 ;
        RECT 7.755 -2.815 8.075 2.535 ;
        RECT 7.755 -12.815 8.075 -7.465 ;
    END
  END RE_BL0
  PIN BL0
    ANTENNADIFFAREA 4.444800 ;
    PORT
      LAYER li1 ;
        RECT 8.300 -2.820 8.470 2.530 ;
        RECT 9.415 0.530 10.755 0.780 ;
        RECT 8.300 -12.820 8.470 -7.470 ;
        RECT 9.415 -9.470 10.755 -9.220 ;
      LAYER mcon ;
        RECT 8.300 2.140 8.470 2.310 ;
        RECT 8.300 1.780 8.470 1.950 ;
        RECT 8.300 1.420 8.470 1.590 ;
        RECT 8.300 1.060 8.470 1.230 ;
        RECT 8.300 0.700 8.470 0.870 ;
        RECT 9.725 0.570 9.895 0.740 ;
        RECT 8.300 0.340 8.470 0.510 ;
        RECT 8.300 -0.020 8.470 0.150 ;
        RECT 8.300 -0.380 8.470 -0.210 ;
        RECT 8.300 -0.740 8.470 -0.570 ;
        RECT 8.300 -1.100 8.470 -0.930 ;
        RECT 8.300 -1.460 8.470 -1.290 ;
        RECT 8.300 -1.820 8.470 -1.650 ;
        RECT 8.300 -2.180 8.470 -2.010 ;
        RECT 8.300 -2.540 8.470 -2.370 ;
        RECT 8.300 -7.860 8.470 -7.690 ;
        RECT 8.300 -8.220 8.470 -8.050 ;
        RECT 8.300 -8.580 8.470 -8.410 ;
        RECT 8.300 -8.940 8.470 -8.770 ;
        RECT 8.300 -9.300 8.470 -9.130 ;
        RECT 9.725 -9.430 9.895 -9.260 ;
        RECT 8.300 -9.660 8.470 -9.490 ;
        RECT 8.300 -10.020 8.470 -9.850 ;
        RECT 8.300 -10.380 8.470 -10.210 ;
        RECT 8.300 -10.740 8.470 -10.570 ;
        RECT 8.300 -11.100 8.470 -10.930 ;
        RECT 8.300 -11.460 8.470 -11.290 ;
        RECT 8.300 -11.820 8.470 -11.650 ;
        RECT 8.300 -12.180 8.470 -12.010 ;
        RECT 8.300 -12.540 8.470 -12.370 ;
      LAYER met1 ;
        RECT 7.960 3.130 8.280 3.390 ;
        RECT 8.060 2.815 8.220 3.130 ;
        RECT 9.105 2.845 9.945 3.405 ;
        RECT 8.060 2.675 8.455 2.815 ;
        RECT 8.315 2.510 8.455 2.675 ;
        RECT 8.270 -2.820 8.500 2.510 ;
        RECT 9.685 0.780 9.945 2.845 ;
        RECT 9.665 0.510 9.955 0.780 ;
        RECT 6.135 -4.200 6.410 -3.980 ;
        RECT 9.685 -4.200 9.945 0.510 ;
        RECT 6.135 -4.405 9.945 -4.200 ;
        RECT 7.960 -6.870 8.280 -6.610 ;
        RECT 8.060 -7.185 8.220 -6.870 ;
        RECT 9.105 -7.155 9.945 -6.595 ;
        RECT 8.060 -7.325 8.455 -7.185 ;
        RECT 8.315 -7.490 8.455 -7.325 ;
        RECT 8.270 -12.820 8.500 -7.490 ;
        RECT 9.685 -9.220 9.945 -7.155 ;
        RECT 9.665 -9.490 9.955 -9.220 ;
        RECT 6.135 -14.200 6.410 -13.980 ;
        RECT 9.685 -14.200 9.945 -9.490 ;
        RECT 6.135 -14.405 9.945 -14.200 ;
      LAYER via ;
        RECT 7.990 3.130 8.250 3.390 ;
        RECT 9.265 3.000 9.525 3.260 ;
        RECT 6.140 -4.350 6.400 -4.090 ;
        RECT 7.990 -6.870 8.250 -6.610 ;
        RECT 9.265 -7.000 9.525 -6.740 ;
        RECT 6.140 -14.350 6.400 -14.090 ;
      LAYER met2 ;
        RECT 4.605 5.570 6.420 7.350 ;
        RECT 6.130 -16.000 6.420 5.570 ;
        RECT 7.990 3.400 8.250 3.420 ;
        RECT 9.105 3.400 9.675 3.410 ;
        RECT 7.990 3.120 9.675 3.400 ;
        RECT 7.990 3.100 8.250 3.120 ;
        RECT 9.105 2.835 9.675 3.120 ;
        RECT 7.990 -6.600 8.250 -6.580 ;
        RECT 9.105 -6.600 9.675 -6.590 ;
        RECT 7.990 -6.880 9.675 -6.600 ;
        RECT 7.990 -6.900 8.250 -6.880 ;
        RECT 9.105 -7.165 9.675 -6.880 ;
    END
  END BL0
  PIN GND
    ANTENNADIFFAREA 0.935600 ;
    PORT
      LAYER li1 ;
        RECT -0.895 3.565 3.010 4.025 ;
        RECT -0.895 -1.395 -0.065 3.565 ;
        RECT 10.765 -0.580 11.015 -0.250 ;
        RECT 20.765 -0.580 21.015 -0.250 ;
        RECT -0.895 -2.230 3.095 -1.395 ;
        RECT 10.740 -2.505 11.000 -1.925 ;
        RECT 20.740 -2.505 21.000 -1.925 ;
        RECT 10.765 -10.580 11.015 -10.250 ;
        RECT 20.765 -10.580 21.015 -10.250 ;
        RECT 10.740 -12.505 11.000 -11.925 ;
        RECT 20.740 -12.505 21.000 -11.925 ;
      LAYER mcon ;
        RECT -0.210 3.720 -0.040 3.890 ;
        RECT 0.260 3.715 0.430 3.885 ;
        RECT 0.785 3.705 0.955 3.875 ;
        RECT 1.255 3.700 1.425 3.870 ;
        RECT 1.680 3.710 1.850 3.880 ;
        RECT 2.150 3.705 2.320 3.875 ;
        RECT 2.675 3.695 2.845 3.865 ;
        RECT -0.590 3.390 -0.420 3.560 ;
        RECT -0.590 2.920 -0.420 3.090 ;
        RECT -0.600 2.385 -0.430 2.555 ;
        RECT -0.595 1.870 -0.425 2.040 ;
        RECT -0.595 1.130 -0.425 1.300 ;
        RECT -0.585 0.590 -0.415 0.760 ;
        RECT -0.595 -0.005 -0.425 0.165 ;
        RECT -0.595 -0.570 -0.425 -0.400 ;
        RECT 10.765 -0.500 10.935 -0.330 ;
        RECT 20.765 -0.500 20.935 -0.330 ;
        RECT -0.575 -1.230 -0.405 -1.060 ;
        RECT -0.585 -1.825 -0.415 -1.655 ;
        RECT -0.115 -1.830 0.055 -1.660 ;
        RECT 0.410 -1.840 0.580 -1.670 ;
        RECT 0.880 -1.845 1.050 -1.675 ;
        RECT 1.305 -1.835 1.475 -1.665 ;
        RECT 1.775 -1.840 1.945 -1.670 ;
        RECT 2.300 -1.850 2.470 -1.680 ;
        RECT 10.790 -2.360 10.960 -2.190 ;
        RECT 20.790 -2.360 20.960 -2.190 ;
        RECT 10.765 -10.500 10.935 -10.330 ;
        RECT 20.765 -10.500 20.935 -10.330 ;
        RECT 10.790 -12.360 10.960 -12.190 ;
        RECT 20.790 -12.360 20.960 -12.190 ;
      LAYER met1 ;
        RECT 8.820 6.285 9.950 7.125 ;
        RECT 2.645 6.060 9.950 6.285 ;
        RECT 2.645 3.965 2.920 6.060 ;
        RECT -0.700 3.625 2.920 3.965 ;
        RECT -0.700 -1.595 -0.310 3.625 ;
        RECT 10.735 -0.260 10.995 0.780 ;
        RECT 20.735 -0.260 20.995 0.780 ;
        RECT 10.675 -0.580 10.995 -0.260 ;
        RECT 20.675 -0.580 20.995 -0.260 ;
        RECT -0.700 -1.960 2.895 -1.595 ;
        RECT 10.735 -3.855 10.995 -0.580 ;
        RECT 13.270 -3.855 13.630 -3.685 ;
        RECT 10.735 -4.060 13.630 -3.855 ;
        RECT 20.735 -3.855 20.995 -0.580 ;
        RECT 23.270 -3.855 23.630 -3.685 ;
        RECT 20.735 -4.060 23.630 -3.855 ;
        RECT 10.735 -10.260 10.995 -9.220 ;
        RECT 20.735 -10.260 20.995 -9.220 ;
        RECT 10.675 -10.580 10.995 -10.260 ;
        RECT 20.675 -10.580 20.995 -10.260 ;
        RECT 10.735 -13.855 10.995 -10.580 ;
        RECT 13.270 -13.855 13.630 -13.685 ;
        RECT 10.735 -14.060 13.630 -13.855 ;
        RECT 20.735 -13.855 20.995 -10.580 ;
        RECT 23.270 -13.855 23.630 -13.685 ;
        RECT 20.735 -14.060 23.630 -13.855 ;
        RECT 13.270 -16.000 24.940 -15.655 ;
      LAYER via ;
        RECT 8.960 6.705 9.220 6.965 ;
        RECT 9.500 6.705 9.760 6.965 ;
        RECT 8.965 6.210 9.225 6.470 ;
        RECT 9.500 6.205 9.760 6.465 ;
        RECT 10.705 -0.550 10.965 -0.290 ;
        RECT 20.705 -0.550 20.965 -0.290 ;
        RECT 13.315 -3.995 13.575 -3.735 ;
        RECT 23.315 -3.995 23.575 -3.735 ;
        RECT 10.705 -10.550 10.965 -10.290 ;
        RECT 20.705 -10.550 20.965 -10.290 ;
        RECT 13.315 -13.995 13.575 -13.735 ;
        RECT 23.315 -13.995 23.575 -13.735 ;
        RECT 13.310 -15.970 13.570 -15.710 ;
        RECT 23.320 -15.965 23.580 -15.705 ;
      LAYER met2 ;
        RECT 8.515 5.570 10.330 7.350 ;
        RECT 10.000 4.265 10.330 5.570 ;
        RECT 10.000 3.920 13.635 4.265 ;
        RECT 9.145 -0.580 11.015 -0.260 ;
        RECT 9.145 -10.580 11.015 -10.260 ;
        RECT 13.270 -16.000 13.635 3.920 ;
        RECT 19.145 -0.580 21.015 -0.260 ;
        RECT 23.265 -3.680 23.630 3.570 ;
        RECT 19.145 -10.580 21.015 -10.260 ;
        RECT 23.270 -16.000 23.635 -3.680 ;
    END
  END GND
  PIN BR0
    ANTENNADIFFAREA 4.444800 ;
    PORT
      LAYER li1 ;
        RECT 9.415 -1.620 10.755 -1.370 ;
        RECT 12.575 -2.820 12.745 2.530 ;
        RECT 9.415 -11.620 10.755 -11.370 ;
        RECT 12.575 -12.820 12.745 -7.470 ;
      LAYER mcon ;
        RECT 12.575 2.140 12.745 2.310 ;
        RECT 12.575 1.780 12.745 1.950 ;
        RECT 12.575 1.420 12.745 1.590 ;
        RECT 12.575 1.060 12.745 1.230 ;
        RECT 12.575 0.700 12.745 0.870 ;
        RECT 12.575 0.340 12.745 0.510 ;
        RECT 12.575 -0.020 12.745 0.150 ;
        RECT 12.575 -0.380 12.745 -0.210 ;
        RECT 12.575 -0.740 12.745 -0.570 ;
        RECT 12.575 -1.100 12.745 -0.930 ;
        RECT 10.265 -1.580 10.435 -1.410 ;
        RECT 12.575 -1.460 12.745 -1.290 ;
        RECT 12.575 -1.820 12.745 -1.650 ;
        RECT 12.575 -2.180 12.745 -2.010 ;
        RECT 12.575 -2.540 12.745 -2.370 ;
        RECT 12.575 -7.860 12.745 -7.690 ;
        RECT 12.575 -8.220 12.745 -8.050 ;
        RECT 12.575 -8.580 12.745 -8.410 ;
        RECT 12.575 -8.940 12.745 -8.770 ;
        RECT 12.575 -9.300 12.745 -9.130 ;
        RECT 12.575 -9.660 12.745 -9.490 ;
        RECT 12.575 -10.020 12.745 -9.850 ;
        RECT 12.575 -10.380 12.745 -10.210 ;
        RECT 12.575 -10.740 12.745 -10.570 ;
        RECT 12.575 -11.100 12.745 -10.930 ;
        RECT 10.265 -11.580 10.435 -11.410 ;
        RECT 12.575 -11.460 12.745 -11.290 ;
        RECT 12.575 -11.820 12.745 -11.650 ;
        RECT 12.575 -12.180 12.745 -12.010 ;
        RECT 12.575 -12.540 12.745 -12.370 ;
      LAYER met1 ;
        RECT 10.205 2.840 11.095 3.420 ;
        RECT 12.235 3.130 12.555 3.390 ;
        RECT 10.205 0.780 10.495 2.840 ;
        RECT 12.335 2.815 12.495 3.130 ;
        RECT 12.335 2.675 12.730 2.815 ;
        RECT 12.590 2.510 12.730 2.675 ;
        RECT 10.215 -1.350 10.475 0.780 ;
        RECT 10.205 -1.620 10.495 -1.350 ;
        RECT 10.215 -4.200 10.475 -1.620 ;
        RECT 12.545 -2.820 12.775 2.510 ;
        RECT 13.910 -4.200 14.185 -3.980 ;
        RECT 10.215 -4.405 14.185 -4.200 ;
        RECT 10.215 -4.410 10.475 -4.405 ;
        RECT 10.205 -7.160 11.095 -6.580 ;
        RECT 12.235 -6.870 12.555 -6.610 ;
        RECT 10.205 -9.220 10.495 -7.160 ;
        RECT 12.335 -7.185 12.495 -6.870 ;
        RECT 12.335 -7.325 12.730 -7.185 ;
        RECT 12.590 -7.490 12.730 -7.325 ;
        RECT 10.215 -11.350 10.475 -9.220 ;
        RECT 10.205 -11.620 10.495 -11.350 ;
        RECT 10.215 -14.200 10.475 -11.620 ;
        RECT 12.545 -12.820 12.775 -7.490 ;
        RECT 13.910 -14.200 14.185 -13.980 ;
        RECT 10.215 -14.405 14.185 -14.200 ;
        RECT 10.215 -14.410 10.475 -14.405 ;
      LAYER via ;
        RECT 10.675 2.990 10.935 3.250 ;
        RECT 12.265 3.130 12.525 3.390 ;
        RECT 13.915 -4.350 14.175 -4.090 ;
        RECT 10.675 -7.010 10.935 -6.750 ;
        RECT 12.265 -6.870 12.525 -6.610 ;
        RECT 13.915 -14.350 14.175 -14.090 ;
      LAYER met2 ;
        RECT 10.470 5.570 12.285 7.350 ;
        RECT 11.975 4.700 12.285 5.570 ;
        RECT 11.975 4.515 14.195 4.700 ;
        RECT 10.500 3.150 12.525 3.420 ;
        RECT 10.500 2.845 11.090 3.150 ;
        RECT 12.265 3.100 12.525 3.150 ;
        RECT 10.500 -6.850 12.525 -6.580 ;
        RECT 10.500 -7.155 11.090 -6.850 ;
        RECT 12.265 -6.900 12.525 -6.850 ;
        RECT 13.905 -16.000 14.195 4.515 ;
    END
  END BR0
  PIN RE_BL1
    ANTENNADIFFAREA 4.200000 ;
    PORT
      LAYER li1 ;
        RECT 17.800 -2.820 17.970 2.530 ;
        RECT 17.800 -12.820 17.970 -7.470 ;
      LAYER mcon ;
        RECT 17.800 2.145 17.970 2.315 ;
        RECT 17.800 1.785 17.970 1.955 ;
        RECT 17.800 1.425 17.970 1.595 ;
        RECT 17.800 1.065 17.970 1.235 ;
        RECT 17.800 0.705 17.970 0.875 ;
        RECT 17.800 0.345 17.970 0.515 ;
        RECT 17.800 -0.015 17.970 0.155 ;
        RECT 17.800 -0.375 17.970 -0.205 ;
        RECT 17.800 -0.735 17.970 -0.565 ;
        RECT 17.800 -1.095 17.970 -0.925 ;
        RECT 17.800 -1.455 17.970 -1.285 ;
        RECT 17.800 -1.815 17.970 -1.645 ;
        RECT 17.800 -2.175 17.970 -2.005 ;
        RECT 17.800 -2.535 17.970 -2.365 ;
        RECT 17.800 -7.855 17.970 -7.685 ;
        RECT 17.800 -8.215 17.970 -8.045 ;
        RECT 17.800 -8.575 17.970 -8.405 ;
        RECT 17.800 -8.935 17.970 -8.765 ;
        RECT 17.800 -9.295 17.970 -9.125 ;
        RECT 17.800 -9.655 17.970 -9.485 ;
        RECT 17.800 -10.015 17.970 -9.845 ;
        RECT 17.800 -10.375 17.970 -10.205 ;
        RECT 17.800 -10.735 17.970 -10.565 ;
        RECT 17.800 -11.095 17.970 -10.925 ;
        RECT 17.800 -11.455 17.970 -11.285 ;
        RECT 17.800 -11.815 17.970 -11.645 ;
        RECT 17.800 -12.175 17.970 -12.005 ;
        RECT 17.800 -12.535 17.970 -12.365 ;
      LAYER met1 ;
        RECT 17.755 -2.465 18.075 2.535 ;
        RECT 15.495 -2.780 18.075 -2.465 ;
        RECT 15.495 -4.925 15.860 -2.780 ;
        RECT 17.755 -2.820 18.075 -2.780 ;
        RECT 17.755 -12.465 18.075 -7.465 ;
        RECT 15.495 -12.780 18.075 -12.465 ;
        RECT 15.495 -14.925 15.860 -12.780 ;
        RECT 17.755 -12.820 18.075 -12.780 ;
      LAYER via ;
        RECT 17.785 2.070 18.045 2.330 ;
        RECT 17.785 1.750 18.045 2.010 ;
        RECT 17.785 1.430 18.045 1.690 ;
        RECT 17.785 1.110 18.045 1.370 ;
        RECT 17.785 0.790 18.045 1.050 ;
        RECT 17.785 0.470 18.045 0.730 ;
        RECT 17.785 0.150 18.045 0.410 ;
        RECT 17.785 -0.170 18.045 0.090 ;
        RECT 17.785 -0.490 18.045 -0.230 ;
        RECT 17.785 -0.810 18.045 -0.550 ;
        RECT 17.785 -1.130 18.045 -0.870 ;
        RECT 17.785 -1.450 18.045 -1.190 ;
        RECT 17.785 -1.770 18.045 -1.510 ;
        RECT 17.785 -2.090 18.045 -1.830 ;
        RECT 17.785 -2.410 18.045 -2.150 ;
        RECT 17.785 -2.730 18.045 -2.470 ;
        RECT 15.565 -4.910 15.825 -4.650 ;
        RECT 17.785 -7.930 18.045 -7.670 ;
        RECT 17.785 -8.250 18.045 -7.990 ;
        RECT 17.785 -8.570 18.045 -8.310 ;
        RECT 17.785 -8.890 18.045 -8.630 ;
        RECT 17.785 -9.210 18.045 -8.950 ;
        RECT 17.785 -9.530 18.045 -9.270 ;
        RECT 17.785 -9.850 18.045 -9.590 ;
        RECT 17.785 -10.170 18.045 -9.910 ;
        RECT 17.785 -10.490 18.045 -10.230 ;
        RECT 17.785 -10.810 18.045 -10.550 ;
        RECT 17.785 -11.130 18.045 -10.870 ;
        RECT 17.785 -11.450 18.045 -11.190 ;
        RECT 17.785 -11.770 18.045 -11.510 ;
        RECT 17.785 -12.090 18.045 -11.830 ;
        RECT 17.785 -12.410 18.045 -12.150 ;
        RECT 17.785 -12.730 18.045 -12.470 ;
        RECT 15.565 -14.910 15.825 -14.650 ;
      LAYER met2 ;
        RECT 14.380 5.570 16.195 7.350 ;
        RECT 15.480 -4.580 15.985 5.570 ;
        RECT 17.755 -2.815 18.075 2.535 ;
        RECT 15.485 -16.000 15.990 -4.580 ;
        RECT 17.755 -12.815 18.075 -7.465 ;
    END
  END RE_BL1
  PIN BL1
    ANTENNADIFFAREA 4.444800 ;
    PORT
      LAYER li1 ;
        RECT 18.300 -2.820 18.470 2.530 ;
        RECT 19.415 0.530 20.755 0.780 ;
        RECT 18.300 -12.820 18.470 -7.470 ;
        RECT 19.415 -9.470 20.755 -9.220 ;
      LAYER mcon ;
        RECT 18.300 2.140 18.470 2.310 ;
        RECT 18.300 1.780 18.470 1.950 ;
        RECT 18.300 1.420 18.470 1.590 ;
        RECT 18.300 1.060 18.470 1.230 ;
        RECT 18.300 0.700 18.470 0.870 ;
        RECT 19.725 0.570 19.895 0.740 ;
        RECT 18.300 0.340 18.470 0.510 ;
        RECT 18.300 -0.020 18.470 0.150 ;
        RECT 18.300 -0.380 18.470 -0.210 ;
        RECT 18.300 -0.740 18.470 -0.570 ;
        RECT 18.300 -1.100 18.470 -0.930 ;
        RECT 18.300 -1.460 18.470 -1.290 ;
        RECT 18.300 -1.820 18.470 -1.650 ;
        RECT 18.300 -2.180 18.470 -2.010 ;
        RECT 18.300 -2.540 18.470 -2.370 ;
        RECT 18.300 -7.860 18.470 -7.690 ;
        RECT 18.300 -8.220 18.470 -8.050 ;
        RECT 18.300 -8.580 18.470 -8.410 ;
        RECT 18.300 -8.940 18.470 -8.770 ;
        RECT 18.300 -9.300 18.470 -9.130 ;
        RECT 19.725 -9.430 19.895 -9.260 ;
        RECT 18.300 -9.660 18.470 -9.490 ;
        RECT 18.300 -10.020 18.470 -9.850 ;
        RECT 18.300 -10.380 18.470 -10.210 ;
        RECT 18.300 -10.740 18.470 -10.570 ;
        RECT 18.300 -11.100 18.470 -10.930 ;
        RECT 18.300 -11.460 18.470 -11.290 ;
        RECT 18.300 -11.820 18.470 -11.650 ;
        RECT 18.300 -12.180 18.470 -12.010 ;
        RECT 18.300 -12.540 18.470 -12.370 ;
      LAYER met1 ;
        RECT 17.960 3.130 18.280 3.390 ;
        RECT 18.060 2.815 18.220 3.130 ;
        RECT 19.105 2.845 19.945 3.405 ;
        RECT 18.060 2.675 18.455 2.815 ;
        RECT 18.315 2.510 18.455 2.675 ;
        RECT 18.270 -2.820 18.500 2.510 ;
        RECT 19.685 0.780 19.945 2.845 ;
        RECT 19.665 0.510 19.955 0.780 ;
        RECT 16.135 -4.200 16.410 -3.980 ;
        RECT 19.685 -4.200 19.945 0.510 ;
        RECT 16.135 -4.405 19.945 -4.200 ;
        RECT 17.960 -6.870 18.280 -6.610 ;
        RECT 18.060 -7.185 18.220 -6.870 ;
        RECT 19.105 -7.155 19.945 -6.595 ;
        RECT 18.060 -7.325 18.455 -7.185 ;
        RECT 18.315 -7.490 18.455 -7.325 ;
        RECT 18.270 -12.820 18.500 -7.490 ;
        RECT 19.685 -9.220 19.945 -7.155 ;
        RECT 19.665 -9.490 19.955 -9.220 ;
        RECT 16.135 -14.200 16.410 -13.980 ;
        RECT 19.685 -14.200 19.945 -9.490 ;
        RECT 16.135 -14.405 19.945 -14.200 ;
      LAYER via ;
        RECT 17.990 3.130 18.250 3.390 ;
        RECT 19.265 3.000 19.525 3.260 ;
        RECT 16.140 -4.350 16.400 -4.090 ;
        RECT 17.990 -6.870 18.250 -6.610 ;
        RECT 19.265 -7.000 19.525 -6.740 ;
        RECT 16.140 -14.350 16.400 -14.090 ;
      LAYER met2 ;
        RECT 16.335 5.570 18.150 7.350 ;
        RECT 16.335 5.220 16.735 5.570 ;
        RECT 16.125 5.055 16.735 5.220 ;
        RECT 16.125 -3.975 16.415 5.055 ;
        RECT 17.990 3.400 18.250 3.420 ;
        RECT 19.105 3.400 19.675 3.410 ;
        RECT 17.990 3.120 19.675 3.400 ;
        RECT 17.990 3.100 18.250 3.120 ;
        RECT 19.105 2.835 19.675 3.120 ;
        RECT 16.130 -16.000 16.420 -3.975 ;
        RECT 17.990 -6.600 18.250 -6.580 ;
        RECT 19.105 -6.600 19.675 -6.590 ;
        RECT 17.990 -6.880 19.675 -6.600 ;
        RECT 17.990 -6.900 18.250 -6.880 ;
        RECT 19.105 -7.165 19.675 -6.880 ;
    END
  END BL1
  PIN RE_BR1
    ANTENNADIFFAREA 4.200000 ;
    PORT
      LAYER li1 ;
        RECT 22.075 -2.820 22.245 2.530 ;
        RECT 22.075 -12.820 22.245 -7.470 ;
      LAYER mcon ;
        RECT 22.075 2.145 22.245 2.315 ;
        RECT 22.075 1.785 22.245 1.955 ;
        RECT 22.075 1.425 22.245 1.595 ;
        RECT 22.075 1.065 22.245 1.235 ;
        RECT 22.075 0.705 22.245 0.875 ;
        RECT 22.075 0.345 22.245 0.515 ;
        RECT 22.075 -0.015 22.245 0.155 ;
        RECT 22.075 -0.375 22.245 -0.205 ;
        RECT 22.075 -0.735 22.245 -0.565 ;
        RECT 22.075 -1.095 22.245 -0.925 ;
        RECT 22.075 -1.455 22.245 -1.285 ;
        RECT 22.075 -1.815 22.245 -1.645 ;
        RECT 22.075 -2.175 22.245 -2.005 ;
        RECT 22.075 -2.535 22.245 -2.365 ;
        RECT 22.075 -7.855 22.245 -7.685 ;
        RECT 22.075 -8.215 22.245 -8.045 ;
        RECT 22.075 -8.575 22.245 -8.405 ;
        RECT 22.075 -8.935 22.245 -8.765 ;
        RECT 22.075 -9.295 22.245 -9.125 ;
        RECT 22.075 -9.655 22.245 -9.485 ;
        RECT 22.075 -10.015 22.245 -9.845 ;
        RECT 22.075 -10.375 22.245 -10.205 ;
        RECT 22.075 -10.735 22.245 -10.565 ;
        RECT 22.075 -11.095 22.245 -10.925 ;
        RECT 22.075 -11.455 22.245 -11.285 ;
        RECT 22.075 -11.815 22.245 -11.645 ;
        RECT 22.075 -12.175 22.245 -12.005 ;
        RECT 22.075 -12.535 22.245 -12.365 ;
      LAYER met1 ;
        RECT 22.030 -3.080 22.350 2.535 ;
        RECT 22.030 -3.285 24.945 -3.080 ;
        RECT 24.665 -4.970 24.945 -3.285 ;
        RECT 22.030 -13.080 22.350 -7.465 ;
        RECT 22.030 -13.285 24.945 -13.080 ;
        RECT 24.665 -14.970 24.945 -13.285 ;
      LAYER via ;
        RECT 22.060 2.070 22.320 2.330 ;
        RECT 22.060 1.750 22.320 2.010 ;
        RECT 22.060 1.430 22.320 1.690 ;
        RECT 22.060 1.110 22.320 1.370 ;
        RECT 22.060 0.790 22.320 1.050 ;
        RECT 22.060 0.470 22.320 0.730 ;
        RECT 22.060 0.150 22.320 0.410 ;
        RECT 22.060 -0.170 22.320 0.090 ;
        RECT 22.060 -0.490 22.320 -0.230 ;
        RECT 22.060 -0.810 22.320 -0.550 ;
        RECT 22.060 -1.130 22.320 -0.870 ;
        RECT 22.060 -1.450 22.320 -1.190 ;
        RECT 22.060 -1.770 22.320 -1.510 ;
        RECT 22.060 -2.090 22.320 -1.830 ;
        RECT 22.060 -2.410 22.320 -2.150 ;
        RECT 22.060 -2.730 22.320 -2.470 ;
        RECT 24.670 -4.910 24.930 -4.650 ;
        RECT 22.060 -7.930 22.320 -7.670 ;
        RECT 22.060 -8.250 22.320 -7.990 ;
        RECT 22.060 -8.570 22.320 -8.310 ;
        RECT 22.060 -8.890 22.320 -8.630 ;
        RECT 22.060 -9.210 22.320 -8.950 ;
        RECT 22.060 -9.530 22.320 -9.270 ;
        RECT 22.060 -9.850 22.320 -9.590 ;
        RECT 22.060 -10.170 22.320 -9.910 ;
        RECT 22.060 -10.490 22.320 -10.230 ;
        RECT 22.060 -10.810 22.320 -10.550 ;
        RECT 22.060 -11.130 22.320 -10.870 ;
        RECT 22.060 -11.450 22.320 -11.190 ;
        RECT 22.060 -11.770 22.320 -11.510 ;
        RECT 22.060 -12.090 22.320 -11.830 ;
        RECT 22.060 -12.410 22.320 -12.150 ;
        RECT 22.060 -12.730 22.320 -12.470 ;
        RECT 24.670 -14.910 24.930 -14.650 ;
      LAYER met2 ;
        RECT 20.245 5.570 22.060 7.350 ;
        RECT 21.795 4.395 22.060 5.570 ;
        RECT 21.795 4.210 24.945 4.395 ;
        RECT 22.030 -2.815 22.350 2.535 ;
        RECT 22.030 -12.815 22.350 -7.465 ;
        RECT 24.440 -14.970 24.945 4.210 ;
        RECT 24.435 -16.000 24.940 -14.970 ;
    END
  END RE_BR1
  PIN BR1
    ANTENNADIFFAREA 4.444800 ;
    PORT
      LAYER li1 ;
        RECT 19.415 -1.620 20.755 -1.370 ;
        RECT 22.575 -2.820 22.745 2.530 ;
        RECT 19.415 -11.620 20.755 -11.370 ;
        RECT 22.575 -12.820 22.745 -7.470 ;
      LAYER mcon ;
        RECT 22.575 2.140 22.745 2.310 ;
        RECT 22.575 1.780 22.745 1.950 ;
        RECT 22.575 1.420 22.745 1.590 ;
        RECT 22.575 1.060 22.745 1.230 ;
        RECT 22.575 0.700 22.745 0.870 ;
        RECT 22.575 0.340 22.745 0.510 ;
        RECT 22.575 -0.020 22.745 0.150 ;
        RECT 22.575 -0.380 22.745 -0.210 ;
        RECT 22.575 -0.740 22.745 -0.570 ;
        RECT 22.575 -1.100 22.745 -0.930 ;
        RECT 20.265 -1.580 20.435 -1.410 ;
        RECT 22.575 -1.460 22.745 -1.290 ;
        RECT 22.575 -1.820 22.745 -1.650 ;
        RECT 22.575 -2.180 22.745 -2.010 ;
        RECT 22.575 -2.540 22.745 -2.370 ;
        RECT 22.575 -7.860 22.745 -7.690 ;
        RECT 22.575 -8.220 22.745 -8.050 ;
        RECT 22.575 -8.580 22.745 -8.410 ;
        RECT 22.575 -8.940 22.745 -8.770 ;
        RECT 22.575 -9.300 22.745 -9.130 ;
        RECT 22.575 -9.660 22.745 -9.490 ;
        RECT 22.575 -10.020 22.745 -9.850 ;
        RECT 22.575 -10.380 22.745 -10.210 ;
        RECT 22.575 -10.740 22.745 -10.570 ;
        RECT 22.575 -11.100 22.745 -10.930 ;
        RECT 20.265 -11.580 20.435 -11.410 ;
        RECT 22.575 -11.460 22.745 -11.290 ;
        RECT 22.575 -11.820 22.745 -11.650 ;
        RECT 22.575 -12.180 22.745 -12.010 ;
        RECT 22.575 -12.540 22.745 -12.370 ;
      LAYER met1 ;
        RECT 20.205 2.840 21.095 3.420 ;
        RECT 22.235 3.130 22.555 3.390 ;
        RECT 20.205 0.780 20.495 2.840 ;
        RECT 22.335 2.815 22.495 3.130 ;
        RECT 22.335 2.675 22.730 2.815 ;
        RECT 22.590 2.510 22.730 2.675 ;
        RECT 20.215 -1.350 20.475 0.780 ;
        RECT 20.205 -1.620 20.495 -1.350 ;
        RECT 20.215 -4.200 20.475 -1.620 ;
        RECT 22.545 -2.820 22.775 2.510 ;
        RECT 23.910 -4.200 24.185 -3.980 ;
        RECT 20.215 -4.405 24.185 -4.200 ;
        RECT 20.215 -4.410 20.475 -4.405 ;
        RECT 20.205 -7.160 21.095 -6.580 ;
        RECT 22.235 -6.870 22.555 -6.610 ;
        RECT 20.205 -9.220 20.495 -7.160 ;
        RECT 22.335 -7.185 22.495 -6.870 ;
        RECT 22.335 -7.325 22.730 -7.185 ;
        RECT 22.590 -7.490 22.730 -7.325 ;
        RECT 20.215 -11.350 20.475 -9.220 ;
        RECT 20.205 -11.620 20.495 -11.350 ;
        RECT 20.215 -14.200 20.475 -11.620 ;
        RECT 22.545 -12.820 22.775 -7.490 ;
        RECT 23.910 -14.200 24.185 -13.980 ;
        RECT 20.215 -14.405 24.185 -14.200 ;
        RECT 20.215 -14.410 20.475 -14.405 ;
      LAYER via ;
        RECT 20.675 2.990 20.935 3.250 ;
        RECT 22.265 3.130 22.525 3.390 ;
        RECT 23.915 -4.350 24.175 -4.090 ;
        RECT 20.675 -7.010 20.935 -6.750 ;
        RECT 22.265 -6.870 22.525 -6.610 ;
        RECT 23.915 -14.350 24.175 -14.090 ;
      LAYER met2 ;
        RECT 18.290 5.570 20.105 7.350 ;
        RECT 19.890 4.070 20.105 5.570 ;
        RECT 19.890 3.925 24.190 4.070 ;
        RECT 20.500 3.150 22.525 3.420 ;
        RECT 20.500 2.845 21.090 3.150 ;
        RECT 22.265 3.100 22.525 3.150 ;
        RECT 23.900 -3.975 24.190 3.925 ;
        RECT 20.500 -6.850 22.525 -6.580 ;
        RECT 20.500 -7.155 21.090 -6.850 ;
        RECT 22.265 -6.900 22.525 -6.850 ;
        RECT 23.905 -16.000 24.195 -3.975 ;
    END
  END BR1
  OBS
      LAYER pwell ;
        RECT 0.390 1.875 1.400 2.495 ;
        RECT 1.605 1.235 2.615 2.495 ;
        RECT 2.660 -0.765 3.670 2.495 ;
        RECT 3.695 -4.775 4.705 2.485 ;
        RECT 7.630 -4.595 8.640 2.665 ;
      LAYER nwell ;
        RECT 8.965 -2.505 9.945 0.780 ;
      LAYER pwell ;
        RECT 10.265 0.340 10.885 0.910 ;
        RECT 10.235 -0.160 10.915 0.340 ;
        RECT 10.235 -0.670 11.145 -0.160 ;
        RECT 10.235 -1.180 10.915 -0.670 ;
        RECT 10.265 -1.750 10.885 -1.180 ;
        RECT 11.905 -4.595 12.915 2.665 ;
        RECT 17.630 -4.595 18.640 2.665 ;
      LAYER nwell ;
        RECT 18.965 -2.505 19.945 0.780 ;
      LAYER pwell ;
        RECT 20.265 0.340 20.885 0.910 ;
        RECT 20.235 -0.160 20.915 0.340 ;
        RECT 20.235 -0.670 21.145 -0.160 ;
        RECT 20.235 -1.180 20.915 -0.670 ;
        RECT 20.265 -1.750 20.885 -1.180 ;
        RECT 21.905 -4.595 22.915 2.665 ;
        RECT 7.630 -14.595 8.640 -7.335 ;
      LAYER nwell ;
        RECT 8.965 -12.505 9.945 -9.220 ;
      LAYER pwell ;
        RECT 10.265 -9.660 10.885 -9.090 ;
        RECT 10.235 -10.160 10.915 -9.660 ;
        RECT 10.235 -10.670 11.145 -10.160 ;
        RECT 10.235 -11.180 10.915 -10.670 ;
        RECT 10.265 -11.750 10.885 -11.180 ;
        RECT 11.905 -14.595 12.915 -7.335 ;
        RECT 17.630 -14.595 18.640 -7.335 ;
      LAYER nwell ;
        RECT 18.965 -12.505 19.945 -9.220 ;
      LAYER pwell ;
        RECT 20.265 -9.660 20.885 -9.090 ;
        RECT 20.235 -10.160 20.915 -9.660 ;
        RECT 20.235 -10.670 21.145 -10.160 ;
        RECT 20.235 -11.180 20.915 -10.670 ;
        RECT 20.265 -11.750 20.885 -11.180 ;
        RECT 21.905 -14.595 22.915 -7.335 ;
      LAYER li1 ;
        RECT 9.425 0.250 10.675 0.360 ;
        RECT 19.425 0.250 20.675 0.360 ;
        RECT 9.345 0.190 10.755 0.250 ;
        RECT 9.345 -0.080 9.745 0.190 ;
        RECT 9.575 -0.410 9.745 -0.080 ;
        RECT 9.925 -0.060 10.255 0.020 ;
        RECT 9.925 -0.230 10.335 -0.060 ;
        RECT 10.505 -0.080 10.755 0.190 ;
        RECT 19.345 0.190 20.755 0.250 ;
        RECT 19.345 -0.080 19.745 0.190 ;
        RECT 10.165 -0.250 10.335 -0.230 ;
        RECT 9.575 -0.580 9.935 -0.410 ;
        RECT 10.165 -0.420 10.595 -0.250 ;
        RECT 9.765 -0.610 9.935 -0.580 ;
        RECT 9.345 -1.030 9.595 -0.760 ;
        RECT 9.765 -0.780 10.255 -0.610 ;
        RECT 9.925 -0.860 10.255 -0.780 ;
        RECT 10.425 -0.760 10.595 -0.420 ;
        RECT 19.575 -0.410 19.745 -0.080 ;
        RECT 19.925 -0.060 20.255 0.020 ;
        RECT 19.925 -0.230 20.335 -0.060 ;
        RECT 20.505 -0.080 20.755 0.190 ;
        RECT 20.165 -0.250 20.335 -0.230 ;
        RECT 19.575 -0.580 19.935 -0.410 ;
        RECT 20.165 -0.420 20.595 -0.250 ;
        RECT 19.765 -0.610 19.935 -0.580 ;
        RECT 10.425 -1.030 10.755 -0.760 ;
        RECT 9.345 -1.090 10.755 -1.030 ;
        RECT 19.345 -1.030 19.595 -0.760 ;
        RECT 19.765 -0.780 20.255 -0.610 ;
        RECT 19.925 -0.860 20.255 -0.780 ;
        RECT 20.425 -0.760 20.595 -0.420 ;
        RECT 20.425 -1.030 20.755 -0.760 ;
        RECT 19.345 -1.090 20.755 -1.030 ;
        RECT 9.425 -1.200 10.675 -1.090 ;
        RECT 19.425 -1.200 20.675 -1.090 ;
        RECT 9.425 -9.750 10.675 -9.640 ;
        RECT 19.425 -9.750 20.675 -9.640 ;
        RECT 9.345 -9.810 10.755 -9.750 ;
        RECT 9.345 -10.080 9.745 -9.810 ;
        RECT 9.575 -10.410 9.745 -10.080 ;
        RECT 9.925 -10.060 10.255 -9.980 ;
        RECT 9.925 -10.230 10.335 -10.060 ;
        RECT 10.505 -10.080 10.755 -9.810 ;
        RECT 19.345 -9.810 20.755 -9.750 ;
        RECT 19.345 -10.080 19.745 -9.810 ;
        RECT 10.165 -10.250 10.335 -10.230 ;
        RECT 9.575 -10.580 9.935 -10.410 ;
        RECT 10.165 -10.420 10.595 -10.250 ;
        RECT 9.765 -10.610 9.935 -10.580 ;
        RECT 9.345 -11.030 9.595 -10.760 ;
        RECT 9.765 -10.780 10.255 -10.610 ;
        RECT 9.925 -10.860 10.255 -10.780 ;
        RECT 10.425 -10.760 10.595 -10.420 ;
        RECT 19.575 -10.410 19.745 -10.080 ;
        RECT 19.925 -10.060 20.255 -9.980 ;
        RECT 19.925 -10.230 20.335 -10.060 ;
        RECT 20.505 -10.080 20.755 -9.810 ;
        RECT 20.165 -10.250 20.335 -10.230 ;
        RECT 19.575 -10.580 19.935 -10.410 ;
        RECT 20.165 -10.420 20.595 -10.250 ;
        RECT 19.765 -10.610 19.935 -10.580 ;
        RECT 10.425 -11.030 10.755 -10.760 ;
        RECT 9.345 -11.090 10.755 -11.030 ;
        RECT 19.345 -11.030 19.595 -10.760 ;
        RECT 19.765 -10.780 20.255 -10.610 ;
        RECT 19.925 -10.860 20.255 -10.780 ;
        RECT 20.425 -10.760 20.595 -10.420 ;
        RECT 20.425 -11.030 20.755 -10.760 ;
        RECT 19.345 -11.090 20.755 -11.030 ;
        RECT 9.425 -11.200 10.675 -11.090 ;
        RECT 19.425 -11.200 20.675 -11.090 ;
      LAYER met2 ;
        RECT 9.145 -1.200 11.015 -0.880 ;
        RECT 19.145 -1.200 21.015 -0.880 ;
        RECT 9.145 -11.200 11.015 -10.880 ;
        RECT 19.145 -11.200 21.015 -10.880 ;
  END
END rram_test
END LIBRARY


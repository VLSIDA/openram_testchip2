VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sky130_sram_1kbyte_1rw_32x256_8
   CLASS BLOCK ;
   SIZE 481.14 BY 223.42 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  116.28 0.0 116.66 1.06 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  121.72 0.0 122.1 1.06 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  127.84 0.0 128.22 1.06 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  133.28 0.0 133.66 1.06 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  139.4 0.0 139.78 1.06 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  146.2 0.0 146.58 1.06 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  150.96 0.0 151.34 1.06 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  157.08 0.0 157.46 1.06 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  162.52 0.0 162.9 1.06 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  168.64 0.0 169.02 1.06 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  174.08 0.0 174.46 1.06 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  180.2 0.0 180.58 1.06 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  186.32 0.0 186.7 1.06 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  191.76 0.0 192.14 1.06 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  198.56 0.0 198.94 1.06 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  204.0 0.0 204.38 1.06 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  210.12 0.0 210.5 1.06 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  216.24 0.0 216.62 1.06 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  221.0 0.0 221.38 1.06 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  227.8 0.0 228.18 1.06 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  233.24 0.0 233.62 1.06 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  239.36 0.0 239.74 1.06 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  245.48 0.0 245.86 1.06 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  250.92 0.0 251.3 1.06 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  256.36 0.0 256.74 1.06 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  262.48 0.0 262.86 1.06 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  268.6 0.0 268.98 1.06 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  274.04 0.0 274.42 1.06 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  279.48 0.0 279.86 1.06 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  285.6 0.0 285.98 1.06 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  291.04 0.0 291.42 1.06 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  297.84 0.0 298.22 1.06 ;
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  302.6 0.0 302.98 1.06 ;
      END
   END din0[32]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  80.92 0.0 81.3 1.06 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  87.04 0.0 87.42 1.06 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 136.68 1.06 137.06 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 144.84 1.06 145.22 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 149.6 1.06 149.98 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  68.0 222.36 68.38 223.42 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  71.4 222.36 71.78 223.42 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  70.72 222.36 71.1 223.42 ;
      END
   END addr0[7]
   PIN addr0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  70.04 222.36 70.42 223.42 ;
      END
   END addr0[8]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 38.76 1.06 39.14 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 47.6 1.06 47.98 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 40.12 1.06 40.5 ;
      END
   END clk0
   PIN wmask0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  93.16 0.0 93.54 1.06 ;
      END
   END wmask0[0]
   PIN wmask0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  98.6 0.0 98.98 1.06 ;
      END
   END wmask0[1]
   PIN wmask0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  105.4 0.0 105.78 1.06 ;
      END
   END wmask0[2]
   PIN wmask0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  110.84 0.0 111.22 1.06 ;
      END
   END wmask0[3]
   PIN spare_wen0
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  309.4 0.0 309.78 1.06 ;
      END
   END spare_wen0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  148.24 0.0 148.62 1.06 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  157.76 0.0 158.14 1.06 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  165.92 0.0 166.3 1.06 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  176.12 0.0 176.5 1.06 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  187.68 0.0 188.06 1.06 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  195.84 0.0 196.22 1.06 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  206.04 0.0 206.42 1.06 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  215.56 0.0 215.94 1.06 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  225.08 0.0 225.46 1.06 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  235.96 0.0 236.34 1.06 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  246.16 0.0 246.54 1.06 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  257.72 0.0 258.1 1.06 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  265.88 0.0 266.26 1.06 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  276.08 0.0 276.46 1.06 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  286.28 0.0 286.66 1.06 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  295.12 0.0 295.5 1.06 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  304.64 0.0 305.02 1.06 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  316.2 0.0 316.58 1.06 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  325.72 0.0 326.1 1.06 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  335.92 0.0 336.3 1.06 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  346.12 0.0 346.5 1.06 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  356.32 0.0 356.7 1.06 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  365.84 0.0 366.22 1.06 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  376.04 0.0 376.42 1.06 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  384.88 0.0 385.26 1.06 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  395.76 0.0 396.14 1.06 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  405.96 0.0 406.34 1.06 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  416.16 0.0 416.54 1.06 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  480.08 66.64 481.14 67.02 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  480.08 57.8 481.14 58.18 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  480.08 61.2 481.14 61.58 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  480.08 63.24 481.14 63.62 ;
      END
   END dout0[31]
   PIN dout0[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER met3 ;
         RECT  480.08 62.56 481.14 62.94 ;
      END
   END dout0[32]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  3.4 3.4 477.74 5.14 ;
         LAYER met4 ;
         RECT  3.4 3.4 5.14 220.02 ;
         LAYER met4 ;
         RECT  476.0 3.4 477.74 220.02 ;
         LAYER met3 ;
         RECT  3.4 218.28 477.74 220.02 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  479.4 0.0 481.14 223.42 ;
         LAYER met4 ;
         RECT  0.0 0.0 1.74 223.42 ;
         LAYER met3 ;
         RECT  0.0 0.0 481.14 1.74 ;
         LAYER met3 ;
         RECT  0.0 221.68 481.14 223.42 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 480.52 222.8 ;
   LAYER  met2 ;
      RECT  0.62 0.62 480.52 222.8 ;
   LAYER  met3 ;
      RECT  1.66 136.08 480.52 137.66 ;
      RECT  0.62 137.66 1.66 144.24 ;
      RECT  0.62 145.82 1.66 149.0 ;
      RECT  0.62 48.58 1.66 136.08 ;
      RECT  0.62 41.1 1.66 47.0 ;
      RECT  1.66 66.04 479.48 67.62 ;
      RECT  1.66 67.62 479.48 136.08 ;
      RECT  479.48 67.62 480.52 136.08 ;
      RECT  479.48 58.78 480.52 60.6 ;
      RECT  479.48 64.22 480.52 66.04 ;
      RECT  1.66 2.8 2.8 5.74 ;
      RECT  1.66 5.74 2.8 66.04 ;
      RECT  2.8 5.74 478.34 66.04 ;
      RECT  478.34 2.8 479.48 5.74 ;
      RECT  478.34 5.74 479.48 66.04 ;
      RECT  1.66 137.66 2.8 217.68 ;
      RECT  1.66 217.68 2.8 220.62 ;
      RECT  2.8 137.66 478.34 217.68 ;
      RECT  478.34 137.66 480.52 217.68 ;
      RECT  478.34 217.68 480.52 220.62 ;
      RECT  0.62 2.34 1.66 38.16 ;
      RECT  479.48 2.34 480.52 57.2 ;
      RECT  1.66 2.34 2.8 2.8 ;
      RECT  2.8 2.34 478.34 2.8 ;
      RECT  478.34 2.34 479.48 2.8 ;
      RECT  0.62 150.58 1.66 221.08 ;
      RECT  1.66 220.62 2.8 221.08 ;
      RECT  2.8 220.62 478.34 221.08 ;
      RECT  478.34 220.62 480.52 221.08 ;
   LAYER  met4 ;
      RECT  115.68 1.66 117.26 222.8 ;
      RECT  117.26 0.62 121.12 1.66 ;
      RECT  122.7 0.62 127.24 1.66 ;
      RECT  128.82 0.62 132.68 1.66 ;
      RECT  134.26 0.62 138.8 1.66 ;
      RECT  140.38 0.62 145.6 1.66 ;
      RECT  151.94 0.62 156.48 1.66 ;
      RECT  169.62 0.62 173.48 1.66 ;
      RECT  181.18 0.62 185.72 1.66 ;
      RECT  199.54 0.62 203.4 1.66 ;
      RECT  217.22 0.62 220.4 1.66 ;
      RECT  228.78 0.62 232.64 1.66 ;
      RECT  240.34 0.62 244.88 1.66 ;
      RECT  251.9 0.62 255.76 1.66 ;
      RECT  269.58 0.62 273.44 1.66 ;
      RECT  280.46 0.62 285.0 1.66 ;
      RECT  298.82 0.62 302.0 1.66 ;
      RECT  81.9 0.62 86.44 1.66 ;
      RECT  67.4 1.66 68.98 221.76 ;
      RECT  68.98 1.66 115.68 221.76 ;
      RECT  72.38 221.76 115.68 222.8 ;
      RECT  68.98 221.76 69.44 222.8 ;
      RECT  88.02 0.62 92.56 1.66 ;
      RECT  94.14 0.62 98.0 1.66 ;
      RECT  99.58 0.62 104.8 1.66 ;
      RECT  106.38 0.62 110.24 1.66 ;
      RECT  111.82 0.62 115.68 1.66 ;
      RECT  147.18 0.62 147.64 1.66 ;
      RECT  149.22 0.62 150.36 1.66 ;
      RECT  158.74 0.62 161.92 1.66 ;
      RECT  163.5 0.62 165.32 1.66 ;
      RECT  166.9 0.62 168.04 1.66 ;
      RECT  175.06 0.62 175.52 1.66 ;
      RECT  177.1 0.62 179.6 1.66 ;
      RECT  188.66 0.62 191.16 1.66 ;
      RECT  192.74 0.62 195.24 1.66 ;
      RECT  196.82 0.62 197.96 1.66 ;
      RECT  204.98 0.62 205.44 1.66 ;
      RECT  207.02 0.62 209.52 1.66 ;
      RECT  211.1 0.62 214.96 1.66 ;
      RECT  221.98 0.62 224.48 1.66 ;
      RECT  226.06 0.62 227.2 1.66 ;
      RECT  234.22 0.62 235.36 1.66 ;
      RECT  236.94 0.62 238.76 1.66 ;
      RECT  247.14 0.62 250.32 1.66 ;
      RECT  258.7 0.62 261.88 1.66 ;
      RECT  263.46 0.62 265.28 1.66 ;
      RECT  266.86 0.62 268.0 1.66 ;
      RECT  275.02 0.62 275.48 1.66 ;
      RECT  277.06 0.62 278.88 1.66 ;
      RECT  287.26 0.62 290.44 1.66 ;
      RECT  292.02 0.62 294.52 1.66 ;
      RECT  296.1 0.62 297.24 1.66 ;
      RECT  303.58 0.62 304.04 1.66 ;
      RECT  305.62 0.62 308.8 1.66 ;
      RECT  310.38 0.62 315.6 1.66 ;
      RECT  317.18 0.62 325.12 1.66 ;
      RECT  326.7 0.62 335.32 1.66 ;
      RECT  336.9 0.62 345.52 1.66 ;
      RECT  347.1 0.62 355.72 1.66 ;
      RECT  357.3 0.62 365.24 1.66 ;
      RECT  366.82 0.62 375.44 1.66 ;
      RECT  377.02 0.62 384.28 1.66 ;
      RECT  385.86 0.62 395.16 1.66 ;
      RECT  396.74 0.62 405.36 1.66 ;
      RECT  406.94 0.62 415.56 1.66 ;
      RECT  2.8 1.66 5.74 2.8 ;
      RECT  2.8 220.62 5.74 221.76 ;
      RECT  5.74 1.66 67.4 2.8 ;
      RECT  5.74 2.8 67.4 220.62 ;
      RECT  5.74 220.62 67.4 221.76 ;
      RECT  117.26 1.66 475.4 2.8 ;
      RECT  117.26 2.8 475.4 220.62 ;
      RECT  117.26 220.62 475.4 222.8 ;
      RECT  475.4 1.66 478.34 2.8 ;
      RECT  475.4 220.62 478.34 222.8 ;
      RECT  417.14 0.62 478.8 1.66 ;
      RECT  478.34 1.66 478.8 2.8 ;
      RECT  478.34 2.8 478.8 220.62 ;
      RECT  478.34 220.62 478.8 222.8 ;
      RECT  2.34 0.62 80.32 1.66 ;
      RECT  2.34 221.76 67.4 222.8 ;
      RECT  2.34 1.66 2.8 2.8 ;
      RECT  2.34 2.8 2.8 220.62 ;
      RECT  2.34 220.62 2.8 221.76 ;
   END
END    sky130_sram_1kbyte_1rw_32x256_8
END    LIBRARY

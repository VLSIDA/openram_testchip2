VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1429.100 2924.800 1430.300 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2228.650 3517.600 2229.210 3524.800 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1904.810 3517.600 1905.370 3524.800 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1580.970 3517.600 1581.530 3524.800 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 933.290 3517.600 933.850 3524.800 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.450 3517.600 610.010 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.610 3517.600 286.170 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3471.140 2.400 3472.340 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3212.740 2.400 3213.940 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2954.340 2.400 2955.540 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1692.940 2924.800 1694.140 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2695.940 2.400 2697.140 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2437.540 2.400 2438.740 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2179.140 2.400 2180.340 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1920.740 2.400 1921.940 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1662.340 2.400 1663.540 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1403.940 2.400 1405.140 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1145.540 2.400 1146.740 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 887.140 2.400 888.340 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 628.740 2.400 629.940 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1956.780 2924.800 1957.980 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2220.620 2924.800 2221.820 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2484.460 2924.800 2485.660 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2748.300 2924.800 2749.500 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3012.140 2924.800 3013.340 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3275.980 2924.800 3277.180 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2876.330 3517.600 2876.890 3524.800 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2552.490 3517.600 2553.050 3524.800 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 43.940 2924.800 45.140 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2286.580 2924.800 2287.780 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2550.420 2924.800 2551.620 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2814.260 2924.800 2815.460 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.100 2924.800 3079.300 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3341.940 2924.800 3343.140 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2795.370 3517.600 2795.930 3524.800 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2471.530 3517.600 2472.090 3524.800 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2147.690 3517.600 2148.250 3524.800 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1823.850 3517.600 1824.410 3524.800 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.010 3517.600 1500.570 3524.800 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 241.820 2924.800 243.020 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1176.170 3517.600 1176.730 3524.800 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 852.330 3517.600 852.890 3524.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.490 3517.600 529.050 3524.800 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 204.650 3517.600 205.210 3524.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3406.540 2.400 3407.740 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3148.140 2.400 3149.340 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2889.740 2.400 2890.940 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2631.340 2.400 2632.540 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2372.940 2.400 2374.140 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2114.540 2.400 2115.740 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 439.700 2924.800 440.900 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1856.140 2.400 1857.340 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1597.740 2.400 1598.940 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1339.340 2.400 1340.540 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1080.940 2.400 1082.140 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 822.540 2.400 823.740 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 564.140 2.400 565.340 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 370.340 2.400 371.540 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 176.540 2.400 177.740 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 637.580 2924.800 638.780 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 835.460 2924.800 836.660 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1033.340 2924.800 1034.540 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1231.220 2924.800 1232.420 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1495.060 2924.800 1496.260 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1758.900 2924.800 1760.100 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2022.740 2924.800 2023.940 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 175.860 2924.800 177.060 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2418.500 2924.800 2419.700 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2682.340 2924.800 2683.540 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2946.180 2924.800 2947.380 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3210.020 2924.800 3211.220 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3473.860 2924.800 3475.060 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2633.450 3517.600 2634.010 3524.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2309.610 3517.600 2310.170 3524.800 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1985.770 3517.600 1986.330 3524.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1661.930 3517.600 1662.490 3524.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 373.740 2924.800 374.940 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1014.250 3517.600 1014.810 3524.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 690.410 3517.600 690.970 3524.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.570 3517.600 367.130 3524.800 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 42.730 3517.600 43.290 3524.800 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3277.340 2.400 3278.540 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3018.940 2.400 3020.140 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2760.540 2.400 2761.740 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2502.140 2.400 2503.340 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2243.740 2.400 2244.940 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1985.340 2.400 1986.540 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 571.620 2924.800 572.820 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1726.940 2.400 1728.140 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1468.540 2.400 1469.740 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1210.140 2.400 1211.340 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 951.740 2.400 952.940 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 693.340 2.400 694.540 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 434.940 2.400 436.140 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 241.140 2.400 242.340 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 47.340 2.400 48.540 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 769.500 2924.800 770.700 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1165.260 2924.800 1166.460 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1363.140 2924.800 1364.340 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1626.980 2924.800 1628.180 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1890.820 2924.800 1892.020 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2154.660 2924.800 2155.860 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 109.900 2924.800 111.100 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2352.540 2924.800 2353.740 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2616.380 2924.800 2617.580 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2880.220 2924.800 2881.420 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3144.060 2924.800 3145.260 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3407.900 2924.800 3409.100 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2714.410 3517.600 2714.970 3524.800 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2390.570 3517.600 2391.130 3524.800 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2066.730 3517.600 2067.290 3524.800 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1742.890 3517.600 1743.450 3524.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 307.780 2924.800 308.980 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1095.210 3517.600 1095.770 3524.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.370 3517.600 771.930 3524.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.530 3517.600 448.090 3524.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.690 3517.600 124.250 3524.800 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3341.940 2.400 3343.140 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3083.540 2.400 3084.740 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2825.140 2.400 2826.340 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2566.740 2.400 2567.940 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2308.340 2.400 2309.540 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2049.940 2.400 2051.140 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 505.660 2924.800 506.860 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1791.540 2.400 1792.740 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1533.140 2.400 1534.340 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1274.740 2.400 1275.940 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1016.340 2.400 1017.540 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 757.940 2.400 759.140 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 499.540 2.400 500.740 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 305.740 2.400 306.940 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 111.940 2.400 113.140 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 703.540 2924.800 704.740 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 901.420 2924.800 902.620 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1099.300 2924.800 1100.500 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1297.180 2924.800 1298.380 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1561.020 2924.800 1562.220 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1824.860 2924.800 1826.060 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2088.700 2924.800 2089.900 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.970 -4.800 684.530 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2339.970 -4.800 2340.530 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2356.530 -4.800 2357.090 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2373.090 -4.800 2373.650 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2389.650 -4.800 2390.210 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2406.210 -4.800 2406.770 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2439.330 -4.800 2439.890 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2455.890 -4.800 2456.450 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2472.450 -4.800 2473.010 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2489.010 -4.800 2489.570 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 849.570 -4.800 850.130 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2505.570 -4.800 2506.130 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2522.130 -4.800 2522.690 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2538.690 -4.800 2539.250 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2555.250 -4.800 2555.810 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2588.370 -4.800 2588.930 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2604.930 -4.800 2605.490 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2621.490 -4.800 2622.050 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2638.050 -4.800 2638.610 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2654.610 -4.800 2655.170 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 866.130 -4.800 866.690 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2671.170 -4.800 2671.730 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2687.730 -4.800 2688.290 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2704.290 -4.800 2704.850 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2720.850 -4.800 2721.410 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2737.410 -4.800 2737.970 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2753.970 -4.800 2754.530 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2770.530 -4.800 2771.090 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2787.090 -4.800 2787.650 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 899.250 -4.800 899.810 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.810 -4.800 916.370 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.370 -4.800 932.930 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.930 -4.800 949.490 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.490 -4.800 966.050 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 982.050 -4.800 982.610 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.610 -4.800 999.170 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.530 -4.800 701.090 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1015.170 -4.800 1015.730 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1031.730 -4.800 1032.290 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1048.290 -4.800 1048.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1064.850 -4.800 1065.410 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1081.410 -4.800 1081.970 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1097.970 -4.800 1098.530 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1131.090 -4.800 1131.650 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1147.650 -4.800 1148.210 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1164.210 -4.800 1164.770 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.090 -4.800 717.650 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1180.770 -4.800 1181.330 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1197.330 -4.800 1197.890 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1213.890 -4.800 1214.450 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1230.450 -4.800 1231.010 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1247.010 -4.800 1247.570 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1263.570 -4.800 1264.130 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1280.130 -4.800 1280.690 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1296.690 -4.800 1297.250 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1313.250 -4.800 1313.810 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1329.810 -4.800 1330.370 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.650 -4.800 734.210 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.930 -4.800 1363.490 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1379.490 -4.800 1380.050 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1396.050 -4.800 1396.610 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1412.610 -4.800 1413.170 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1429.170 -4.800 1429.730 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1445.730 -4.800 1446.290 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1462.290 -4.800 1462.850 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1478.850 -4.800 1479.410 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 750.210 -4.800 750.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1511.970 -4.800 1512.530 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1528.530 -4.800 1529.090 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1545.090 -4.800 1545.650 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1561.650 -4.800 1562.210 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1578.210 -4.800 1578.770 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1594.770 -4.800 1595.330 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1611.330 -4.800 1611.890 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1627.890 -4.800 1628.450 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1644.450 -4.800 1645.010 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1661.010 -4.800 1661.570 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.770 -4.800 767.330 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1677.570 -4.800 1678.130 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1694.130 -4.800 1694.690 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1710.690 -4.800 1711.250 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1743.810 -4.800 1744.370 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1760.370 -4.800 1760.930 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1776.930 -4.800 1777.490 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1793.490 -4.800 1794.050 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1810.050 -4.800 1810.610 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1826.610 -4.800 1827.170 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 783.330 -4.800 783.890 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1843.170 -4.800 1843.730 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1859.730 -4.800 1860.290 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1876.290 -4.800 1876.850 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1892.850 -4.800 1893.410 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1909.410 -4.800 1909.970 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1925.970 -4.800 1926.530 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1942.530 -4.800 1943.090 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1975.650 -4.800 1976.210 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1992.210 -4.800 1992.770 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 799.890 -4.800 800.450 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2008.770 -4.800 2009.330 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2025.330 -4.800 2025.890 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2041.890 -4.800 2042.450 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2058.450 -4.800 2059.010 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2075.010 -4.800 2075.570 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2091.570 -4.800 2092.130 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2108.130 -4.800 2108.690 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2124.690 -4.800 2125.250 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2141.250 -4.800 2141.810 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2157.810 -4.800 2158.370 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 816.450 -4.800 817.010 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2174.370 -4.800 2174.930 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2207.490 -4.800 2208.050 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2224.050 -4.800 2224.610 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2240.610 -4.800 2241.170 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2257.170 -4.800 2257.730 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2273.730 -4.800 2274.290 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2290.290 -4.800 2290.850 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2306.850 -4.800 2307.410 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2323.410 -4.800 2323.970 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 833.010 -4.800 833.570 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.490 -4.800 690.050 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2362.050 -4.800 2362.610 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2378.610 -4.800 2379.170 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2395.170 -4.800 2395.730 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2411.730 -4.800 2412.290 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2428.290 -4.800 2428.850 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2444.850 -4.800 2445.410 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2461.410 -4.800 2461.970 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2477.970 -4.800 2478.530 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 855.090 -4.800 855.650 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2511.090 -4.800 2511.650 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2527.650 -4.800 2528.210 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2544.210 -4.800 2544.770 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2560.770 -4.800 2561.330 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2577.330 -4.800 2577.890 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2593.890 -4.800 2594.450 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2610.450 -4.800 2611.010 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2627.010 -4.800 2627.570 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2643.570 -4.800 2644.130 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2660.130 -4.800 2660.690 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.650 -4.800 872.210 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2676.690 -4.800 2677.250 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2693.250 -4.800 2693.810 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2709.810 -4.800 2710.370 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2742.930 -4.800 2743.490 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2759.490 -4.800 2760.050 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2776.050 -4.800 2776.610 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2792.610 -4.800 2793.170 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 888.210 -4.800 888.770 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.770 -4.800 905.330 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 921.330 -4.800 921.890 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.890 -4.800 938.450 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 954.450 -4.800 955.010 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 971.010 -4.800 971.570 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 987.570 -4.800 988.130 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1004.130 -4.800 1004.690 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.050 -4.800 706.610 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1020.690 -4.800 1021.250 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.810 -4.800 1054.370 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1070.370 -4.800 1070.930 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1086.930 -4.800 1087.490 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1103.490 -4.800 1104.050 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.050 -4.800 1120.610 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1136.610 -4.800 1137.170 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1153.170 -4.800 1153.730 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1169.730 -4.800 1170.290 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.610 -4.800 723.170 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1186.290 -4.800 1186.850 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.850 -4.800 1203.410 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1219.410 -4.800 1219.970 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1235.970 -4.800 1236.530 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1252.530 -4.800 1253.090 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1285.650 -4.800 1286.210 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1302.210 -4.800 1302.770 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1318.770 -4.800 1319.330 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1335.330 -4.800 1335.890 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.170 -4.800 739.730 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1351.890 -4.800 1352.450 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1368.450 -4.800 1369.010 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1385.010 -4.800 1385.570 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1401.570 -4.800 1402.130 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1434.690 -4.800 1435.250 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1451.250 -4.800 1451.810 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1467.810 -4.800 1468.370 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1484.370 -4.800 1484.930 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.930 -4.800 1501.490 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 755.730 -4.800 756.290 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1517.490 -4.800 1518.050 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1534.050 -4.800 1534.610 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1550.610 -4.800 1551.170 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1567.170 -4.800 1567.730 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1583.730 -4.800 1584.290 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1600.290 -4.800 1600.850 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.850 -4.800 1617.410 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1633.410 -4.800 1633.970 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1666.530 -4.800 1667.090 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.290 -4.800 772.850 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1683.090 -4.800 1683.650 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1699.650 -4.800 1700.210 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1716.210 -4.800 1716.770 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1732.770 -4.800 1733.330 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1749.330 -4.800 1749.890 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1765.890 -4.800 1766.450 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1782.450 -4.800 1783.010 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1799.010 -4.800 1799.570 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1815.570 -4.800 1816.130 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1832.130 -4.800 1832.690 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.850 -4.800 789.410 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1848.690 -4.800 1849.250 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1865.250 -4.800 1865.810 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1898.370 -4.800 1898.930 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1914.930 -4.800 1915.490 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1931.490 -4.800 1932.050 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1948.050 -4.800 1948.610 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1964.610 -4.800 1965.170 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1981.170 -4.800 1981.730 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1997.730 -4.800 1998.290 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2014.290 -4.800 2014.850 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2030.850 -4.800 2031.410 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2047.410 -4.800 2047.970 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2063.970 -4.800 2064.530 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2080.530 -4.800 2081.090 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2097.090 -4.800 2097.650 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2130.210 -4.800 2130.770 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2146.770 -4.800 2147.330 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2163.330 -4.800 2163.890 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.970 -4.800 822.530 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2179.890 -4.800 2180.450 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2196.450 -4.800 2197.010 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2213.010 -4.800 2213.570 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2229.570 -4.800 2230.130 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2246.130 -4.800 2246.690 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2262.690 -4.800 2263.250 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2279.250 -4.800 2279.810 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2295.810 -4.800 2296.370 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2312.370 -4.800 2312.930 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2328.930 -4.800 2329.490 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 838.530 -4.800 839.090 2.400 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.010 -4.800 695.570 2.400 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2351.010 -4.800 2351.570 2.400 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2367.570 -4.800 2368.130 2.400 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2384.130 -4.800 2384.690 2.400 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2400.690 -4.800 2401.250 2.400 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2433.810 -4.800 2434.370 2.400 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2450.370 -4.800 2450.930 2.400 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2466.930 -4.800 2467.490 2.400 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2483.490 -4.800 2484.050 2.400 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2500.050 -4.800 2500.610 2.400 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.610 -4.800 861.170 2.400 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2516.610 -4.800 2517.170 2.400 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2533.170 -4.800 2533.730 2.400 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2549.730 -4.800 2550.290 2.400 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2566.290 -4.800 2566.850 2.400 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2582.850 -4.800 2583.410 2.400 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2599.410 -4.800 2599.970 2.400 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2615.970 -4.800 2616.530 2.400 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2632.530 -4.800 2633.090 2.400 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2665.650 -4.800 2666.210 2.400 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.170 -4.800 877.730 2.400 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2682.210 -4.800 2682.770 2.400 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2698.770 -4.800 2699.330 2.400 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2715.330 -4.800 2715.890 2.400 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2731.890 -4.800 2732.450 2.400 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2748.450 -4.800 2749.010 2.400 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2765.010 -4.800 2765.570 2.400 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2781.570 -4.800 2782.130 2.400 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2798.130 -4.800 2798.690 2.400 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.730 -4.800 894.290 2.400 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 910.290 -4.800 910.850 2.400 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.850 -4.800 927.410 2.400 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 943.410 -4.800 943.970 2.400 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.530 -4.800 977.090 2.400 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 993.090 -4.800 993.650 2.400 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1009.650 -4.800 1010.210 2.400 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.570 -4.800 712.130 2.400 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1026.210 -4.800 1026.770 2.400 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1042.770 -4.800 1043.330 2.400 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1059.330 -4.800 1059.890 2.400 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1075.890 -4.800 1076.450 2.400 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1092.450 -4.800 1093.010 2.400 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1109.010 -4.800 1109.570 2.400 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1125.570 -4.800 1126.130 2.400 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1142.130 -4.800 1142.690 2.400 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1158.690 -4.800 1159.250 2.400 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.250 -4.800 1175.810 2.400 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 728.130 -4.800 728.690 2.400 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.370 -4.800 1208.930 2.400 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1224.930 -4.800 1225.490 2.400 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1241.490 -4.800 1242.050 2.400 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1258.050 -4.800 1258.610 2.400 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1274.610 -4.800 1275.170 2.400 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.170 -4.800 1291.730 2.400 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1307.730 -4.800 1308.290 2.400 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1324.290 -4.800 1324.850 2.400 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1340.850 -4.800 1341.410 2.400 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.690 -4.800 745.250 2.400 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1357.410 -4.800 1357.970 2.400 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1373.970 -4.800 1374.530 2.400 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1390.530 -4.800 1391.090 2.400 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1407.090 -4.800 1407.650 2.400 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1440.210 -4.800 1440.770 2.400 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1456.770 -4.800 1457.330 2.400 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1473.330 -4.800 1473.890 2.400 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1489.890 -4.800 1490.450 2.400 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1506.450 -4.800 1507.010 2.400 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 761.250 -4.800 761.810 2.400 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1523.010 -4.800 1523.570 2.400 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1539.570 -4.800 1540.130 2.400 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1556.130 -4.800 1556.690 2.400 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1589.250 -4.800 1589.810 2.400 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1605.810 -4.800 1606.370 2.400 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1622.370 -4.800 1622.930 2.400 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1638.930 -4.800 1639.490 2.400 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1655.490 -4.800 1656.050 2.400 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1672.050 -4.800 1672.610 2.400 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.810 -4.800 778.370 2.400 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1688.610 -4.800 1689.170 2.400 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1705.170 -4.800 1705.730 2.400 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1721.730 -4.800 1722.290 2.400 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1738.290 -4.800 1738.850 2.400 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1754.850 -4.800 1755.410 2.400 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1771.410 -4.800 1771.970 2.400 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.970 -4.800 1788.530 2.400 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1821.090 -4.800 1821.650 2.400 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1837.650 -4.800 1838.210 2.400 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.370 -4.800 794.930 2.400 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1854.210 -4.800 1854.770 2.400 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1870.770 -4.800 1871.330 2.400 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1887.330 -4.800 1887.890 2.400 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1903.890 -4.800 1904.450 2.400 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1920.450 -4.800 1921.010 2.400 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1937.010 -4.800 1937.570 2.400 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1953.570 -4.800 1954.130 2.400 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1970.130 -4.800 1970.690 2.400 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1986.690 -4.800 1987.250 2.400 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2003.250 -4.800 2003.810 2.400 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.930 -4.800 811.490 2.400 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2019.810 -4.800 2020.370 2.400 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2052.930 -4.800 2053.490 2.400 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2069.490 -4.800 2070.050 2.400 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2086.050 -4.800 2086.610 2.400 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2102.610 -4.800 2103.170 2.400 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2119.170 -4.800 2119.730 2.400 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2135.730 -4.800 2136.290 2.400 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2152.290 -4.800 2152.850 2.400 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2168.850 -4.800 2169.410 2.400 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.490 -4.800 828.050 2.400 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2185.410 -4.800 2185.970 2.400 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2201.970 -4.800 2202.530 2.400 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2218.530 -4.800 2219.090 2.400 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2235.090 -4.800 2235.650 2.400 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2251.650 -4.800 2252.210 2.400 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2284.770 -4.800 2285.330 2.400 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2301.330 -4.800 2301.890 2.400 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2317.890 -4.800 2318.450 2.400 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2334.450 -4.800 2335.010 2.400 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 844.050 -4.800 844.610 2.400 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2809.170 -4.800 2809.730 2.400 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2814.690 -4.800 2815.250 2.400 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2820.210 -4.800 2820.770 2.400 ;
    END
  END user_irq[2]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -11.580 -6.220 -8.480 3525.900 ;
    END
    PORT
      LAYER met5 ;
        RECT -11.580 -6.220 2931.200 -3.120 ;
    END
    PORT
      LAYER met5 ;
        RECT -11.580 3522.800 2931.200 3525.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 2928.100 -6.220 2931.200 3525.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 8.970 -39.820 12.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 -39.820 192.070 167.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 410.420 192.070 567.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 1006.000 192.070 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 2157.140 192.070 2310.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 2734.360 192.070 2885.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 3352.380 192.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 -39.820 372.070 167.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 410.420 372.070 567.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 1006.000 372.070 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 2157.140 372.070 2310.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 2734.360 372.070 2885.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 3352.380 372.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 -39.820 552.070 167.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 410.420 552.070 567.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 1006.000 552.070 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 2157.140 552.070 2310.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 2734.360 552.070 2885.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 3352.380 552.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 -39.820 732.070 567.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 1006.000 732.070 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 2157.140 732.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.970 -39.820 912.070 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.970 2157.140 912.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.970 -39.820 1092.070 990.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.970 1247.250 1092.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1268.970 -39.820 1272.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1448.970 -39.820 1452.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1628.970 -39.820 1632.070 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1628.970 613.620 1632.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.970 -39.820 1812.070 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.970 613.620 1812.070 786.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.970 1224.580 1812.070 1494.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.970 1840.760 1812.070 2050.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.970 2742.900 1812.070 3018.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.970 3365.040 1812.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1988.970 -39.820 1992.070 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1988.970 613.620 1992.070 786.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1988.970 1224.580 1992.070 1494.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 1988.970 1840.760 1992.070 2050.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 1988.970 2742.900 1992.070 3018.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1988.970 3365.040 1992.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 -39.820 2172.070 786.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 1224.580 2172.070 1494.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 1840.760 2172.070 2050.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 2742.900 2172.070 3018.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 3365.040 2172.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.970 -39.820 2352.070 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.970 613.620 2352.070 786.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.970 1224.580 2352.070 2050.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.970 2742.900 2352.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 -39.820 2532.070 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 613.620 2532.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.970 -39.820 2712.070 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.970 613.620 2712.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2888.970 -39.820 2892.070 3559.500 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 14.330 2964.800 17.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 194.330 2964.800 197.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 374.330 2964.800 377.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 554.330 2964.800 557.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 734.330 2964.800 737.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 914.330 2964.800 917.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1094.330 2964.800 1097.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1274.330 2964.800 1277.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1454.330 2964.800 1457.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1634.330 2964.800 1637.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1814.330 2964.800 1817.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1994.330 2964.800 1997.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2174.330 2964.800 2177.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2354.330 2964.800 2357.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2534.330 2964.800 2537.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2714.330 2964.800 2717.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2894.330 2964.800 2897.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3074.330 2964.800 3077.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3254.330 2964.800 3257.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3434.330 2964.800 3437.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 8.970 2771.150 732.070 2774.250 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -21.180 -15.820 -18.080 3535.500 ;
    END
    PORT
      LAYER met5 ;
        RECT -21.180 -15.820 2940.800 -12.720 ;
    END
    PORT
      LAYER met5 ;
        RECT -21.180 3532.400 2940.800 3535.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2937.700 -15.820 2940.800 3535.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 53.970 -39.820 57.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 233.970 -39.820 237.070 167.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 233.970 1006.000 237.070 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 233.970 3352.380 237.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 413.970 -39.820 417.070 167.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 413.970 1006.000 417.070 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 413.970 3352.380 417.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 593.970 -39.820 597.070 167.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 593.970 1006.000 597.070 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 593.970 3352.380 597.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 773.970 -39.820 777.070 567.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 773.970 1006.000 777.070 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 773.970 2157.140 777.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 953.970 -39.820 957.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1133.970 -39.820 1137.070 990.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1133.970 1247.250 1137.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1313.970 -39.820 1317.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1493.970 -39.820 1497.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1673.970 -39.820 1677.070 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1673.970 613.620 1677.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1853.970 -39.820 1857.070 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1853.970 1840.760 1857.070 2050.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 1853.970 2742.900 1857.070 3018.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1853.970 3365.040 1857.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2033.970 -39.820 2037.070 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2033.970 1840.760 2037.070 2050.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 2033.970 2742.900 2037.070 3018.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2033.970 3365.040 2037.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2213.970 -39.820 2217.070 786.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2213.970 1224.580 2217.070 2050.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 2213.970 2742.900 2217.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2393.970 -39.820 2397.070 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2393.970 1224.580 2397.070 2050.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 2393.970 2742.900 2397.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2573.970 -39.820 2577.070 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2573.970 613.620 2577.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2753.970 -39.820 2757.070 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2753.970 613.620 2757.070 3559.500 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 59.330 2964.800 62.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 239.330 2964.800 242.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 419.330 2964.800 422.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 599.330 2964.800 602.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 779.330 2964.800 782.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 959.330 2964.800 962.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1139.330 2964.800 1142.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1319.330 2964.800 1322.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1499.330 2964.800 1502.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1679.330 2964.800 1682.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1859.330 2964.800 1862.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2039.330 2964.800 2042.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2219.330 2964.800 2222.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2399.330 2964.800 2402.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2579.330 2964.800 2582.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2759.330 2964.800 2762.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2939.330 2964.800 2942.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3119.330 2964.800 3122.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3299.330 2964.800 3302.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3479.330 2964.800 3482.430 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -30.780 -25.420 -27.680 3545.100 ;
    END
    PORT
      LAYER met5 ;
        RECT -30.780 -25.420 2950.400 -22.320 ;
    END
    PORT
      LAYER met5 ;
        RECT -30.780 3542.000 2950.400 3545.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 2947.300 -25.420 2950.400 3545.100 ;
    END
    PORT
      LAYER met4 ;
        RECT 98.970 -39.820 102.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.970 -39.820 282.070 167.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.970 1006.000 282.070 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 -39.820 462.070 167.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 1006.000 462.070 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 -39.820 642.070 167.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 1006.000 642.070 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 818.970 -39.820 822.070 567.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 818.970 1006.000 822.070 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 818.970 2157.140 822.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 998.970 -39.820 1002.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1178.970 -39.820 1182.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1358.970 -39.820 1362.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1538.970 -39.820 1542.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1718.970 -39.820 1722.070 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1718.970 2742.900 1722.070 3018.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1898.970 -39.820 1902.070 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1898.970 2742.900 1902.070 3018.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2078.970 -39.820 2082.070 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2078.970 2742.900 2082.070 3018.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 -39.820 2262.070 786.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 1224.580 2262.070 2050.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 2742.900 2262.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2438.970 -39.820 2442.070 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2438.970 613.620 2442.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2618.970 -39.820 2622.070 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2618.970 613.620 2622.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2798.970 -39.820 2802.070 3559.500 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 104.330 2964.800 107.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 284.330 2964.800 287.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 464.330 2964.800 467.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 644.330 2964.800 647.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 824.330 2964.800 827.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1004.330 2964.800 1007.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1184.330 2964.800 1187.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1364.330 2964.800 1367.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1544.330 2964.800 1547.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1724.330 2964.800 1727.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1904.330 2964.800 1907.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2084.330 2964.800 2087.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2264.330 2964.800 2267.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2444.330 2964.800 2447.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2624.330 2964.800 2627.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2804.330 2964.800 2807.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2984.330 2964.800 2987.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3164.330 2964.800 3167.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3344.330 2964.800 3347.430 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -40.380 -35.020 -37.280 3554.700 ;
    END
    PORT
      LAYER met5 ;
        RECT -40.380 -35.020 2960.000 -31.920 ;
    END
    PORT
      LAYER met5 ;
        RECT -40.380 3551.600 2960.000 3554.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2956.900 -35.020 2960.000 3554.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 143.970 -39.820 147.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 323.970 -39.820 327.070 167.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 323.970 1006.000 327.070 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 323.970 3352.380 327.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 503.970 -39.820 507.070 167.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 503.970 1006.000 507.070 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 503.970 3352.380 507.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 683.970 -39.820 687.070 167.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 683.970 1006.000 687.070 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 683.970 2734.360 687.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 863.970 -39.820 867.070 567.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 863.970 1006.000 867.070 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 863.970 2157.140 867.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1043.970 -39.820 1047.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1223.970 -39.820 1227.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.970 -39.820 1407.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1583.970 -39.820 1587.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1763.970 -39.820 1767.070 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1763.970 1224.580 1767.070 1494.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 1763.970 3365.040 1767.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1943.970 -39.820 1947.070 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1943.970 1224.580 1947.070 1494.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 1943.970 3365.040 1947.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2123.970 -39.820 2127.070 786.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2123.970 1224.580 2127.070 1494.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 2123.970 3365.040 2127.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2303.970 -39.820 2307.070 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2303.970 1224.580 2307.070 2050.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 2303.970 2742.900 2307.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2483.970 -39.820 2487.070 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2483.970 613.620 2487.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2663.970 -39.820 2667.070 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2663.970 613.620 2667.070 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2843.970 -39.820 2847.070 3559.500 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 149.330 2964.800 152.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 329.330 2964.800 332.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 509.330 2964.800 512.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 689.330 2964.800 692.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 869.330 2964.800 872.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1049.330 2964.800 1052.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1229.330 2964.800 1232.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1409.330 2964.800 1412.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1589.330 2964.800 1592.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1769.330 2964.800 1772.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1949.330 2964.800 1952.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2129.330 2964.800 2132.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2309.330 2964.800 2312.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2489.330 2964.800 2492.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2669.330 2964.800 2672.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2849.330 2964.800 2852.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3029.330 2964.800 3032.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3209.330 2964.800 3212.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3389.330 2964.800 3392.430 ;
    END
  END vdda2
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -35.580 -30.220 -32.480 3549.900 ;
    END
    PORT
      LAYER met5 ;
        RECT -35.580 -30.220 2955.200 -27.120 ;
    END
    PORT
      LAYER met5 ;
        RECT -35.580 3546.800 2955.200 3549.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 2952.100 -30.220 2955.200 3549.900 ;
    END
    PORT
      LAYER met4 ;
        RECT 121.470 -39.820 124.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 301.470 -39.820 304.570 167.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 301.470 1006.000 304.570 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 301.470 3352.380 304.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.470 -39.820 484.570 167.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.470 1006.000 484.570 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.470 3352.380 484.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 661.470 -39.820 664.570 167.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 661.470 1006.000 664.570 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 661.470 3352.380 664.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 841.470 -39.820 844.570 567.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 841.470 1006.000 844.570 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 841.470 2157.140 844.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1021.470 -39.820 1024.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1201.470 -39.820 1204.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1381.470 -39.820 1384.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1561.470 -39.820 1564.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1741.470 -39.820 1744.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1741.470 2742.900 1744.570 3018.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1741.470 3365.040 1744.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1921.470 -39.820 1924.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1921.470 2742.900 1924.570 3018.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1921.470 3365.040 1924.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2101.470 -39.820 2104.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2101.470 2742.900 2104.570 3018.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2101.470 3365.040 2104.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2281.470 -39.820 2284.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2281.470 1224.580 2284.570 2050.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 2281.470 2742.900 2284.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2461.470 -39.820 2464.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2461.470 613.620 2464.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2641.470 -39.820 2644.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2641.470 613.620 2644.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2821.470 -39.820 2824.570 3559.500 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 126.830 2964.800 129.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 306.830 2964.800 309.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 486.830 2964.800 489.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 666.830 2964.800 669.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 846.830 2964.800 849.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1026.830 2964.800 1029.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1206.830 2964.800 1209.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1386.830 2964.800 1389.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1566.830 2964.800 1569.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1746.830 2964.800 1749.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1926.830 2964.800 1929.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2106.830 2964.800 2109.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2286.830 2964.800 2289.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2466.830 2964.800 2469.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2646.830 2964.800 2649.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2826.830 2964.800 2829.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3006.830 2964.800 3009.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3186.830 2964.800 3189.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3366.830 2964.800 3369.930 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -45.180 -39.820 -42.080 3559.500 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 -39.820 2964.800 -36.720 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3556.400 2964.800 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2961.700 -39.820 2964.800 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 166.470 -39.820 169.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 346.470 1006.000 349.570 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 346.470 3352.380 349.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 526.470 1006.000 529.570 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 526.470 3352.380 529.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 706.470 -39.820 709.570 567.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 706.470 1006.000 709.570 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 706.470 2157.140 709.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 886.470 -39.820 889.570 567.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 886.470 1006.000 889.570 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 886.470 2157.140 889.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1066.470 -39.820 1069.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1246.470 -39.820 1249.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1426.470 -39.820 1429.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1606.470 -39.820 1609.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1606.470 613.620 1609.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1786.470 -39.820 1789.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1786.470 1224.580 1789.570 1494.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 1786.470 3365.040 1789.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1966.470 -39.820 1969.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1966.470 1224.580 1969.570 1494.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 1966.470 3365.040 1969.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2146.470 -39.820 2149.570 786.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2146.470 1224.580 2149.570 1494.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 2146.470 3365.040 2149.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2326.470 -39.820 2329.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2326.470 1224.580 2329.570 2050.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 2326.470 2742.900 2329.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2506.470 -39.820 2509.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2506.470 613.620 2509.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2686.470 -39.820 2689.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2686.470 613.620 2689.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2866.470 -39.820 2869.570 3559.500 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 171.830 2964.800 174.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 351.830 2964.800 354.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 531.830 2964.800 534.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 711.830 2964.800 714.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 891.830 2964.800 894.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1071.830 2964.800 1074.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1251.830 2964.800 1254.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1431.830 2964.800 1434.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1611.830 2964.800 1614.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1791.830 2964.800 1794.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1971.830 2964.800 1974.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2151.830 2964.800 2154.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2331.830 2964.800 2334.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2511.830 2964.800 2514.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2691.830 2964.800 2694.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2871.830 2964.800 2874.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3051.830 2964.800 3054.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3231.830 2964.800 3234.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3411.830 2964.800 3414.930 ;
    END
  END vssa2
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -16.380 -11.020 -13.280 3530.700 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 -11.020 2936.000 -7.920 ;
    END
    PORT
      LAYER met5 ;
        RECT -16.380 3527.600 2936.000 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 2932.900 -11.020 2936.000 3530.700 ;
    END
    PORT
      LAYER met4 ;
        RECT 31.470 -39.820 34.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 211.470 -39.820 214.570 167.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 211.470 410.420 214.570 567.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 211.470 1006.000 214.570 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 211.470 2157.140 214.570 2310.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 211.470 2734.360 214.570 2885.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 211.470 3352.380 214.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 391.470 -39.820 394.570 167.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 391.470 410.420 394.570 567.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 391.470 1006.000 394.570 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 391.470 2157.140 394.570 2310.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 391.470 2734.360 394.570 2885.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 391.470 3352.380 394.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 571.470 -39.820 574.570 167.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 571.470 410.420 574.570 567.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 571.470 1006.000 574.570 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 571.470 2157.140 574.570 2310.740 ;
    END
    PORT
      LAYER met4 ;
        RECT 571.470 2734.360 574.570 2885.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 571.470 3352.380 574.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 751.470 -39.820 754.570 567.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 751.470 1006.000 754.570 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 751.470 2157.140 754.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 931.470 -39.820 934.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1111.470 -39.820 1114.570 990.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1111.470 1247.250 1114.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1291.470 -39.820 1294.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1471.470 -39.820 1474.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1651.470 -39.820 1654.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1651.470 613.620 1654.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1831.470 -39.820 1834.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1831.470 613.620 1834.570 786.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1831.470 1224.580 1834.570 1494.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 1831.470 1840.760 1834.570 2050.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 1831.470 2742.900 1834.570 3018.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1831.470 3365.040 1834.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2011.470 -39.820 2014.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2011.470 613.620 2014.570 786.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2011.470 1224.580 2014.570 1494.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 2011.470 1840.760 2014.570 2050.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 2011.470 2742.900 2014.570 3018.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2011.470 3365.040 2014.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2191.470 -39.820 2194.570 786.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2191.470 1224.580 2194.570 1494.660 ;
    END
    PORT
      LAYER met4 ;
        RECT 2191.470 1840.760 2194.570 2050.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 2191.470 2742.900 2194.570 3018.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2191.470 3365.040 2194.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2371.470 -39.820 2374.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2371.470 613.620 2374.570 786.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2371.470 1224.580 2374.570 2050.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 2371.470 2742.900 2374.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2551.470 -39.820 2554.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2551.470 613.620 2554.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2731.470 -39.820 2734.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2731.470 613.620 2734.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2911.470 -39.820 2914.570 3559.500 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 36.830 2964.800 39.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 216.830 2964.800 219.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 396.830 2964.800 399.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 576.830 2964.800 579.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 756.830 2964.800 759.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 936.830 2964.800 939.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1116.830 2964.800 1119.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1296.830 2964.800 1299.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1476.830 2964.800 1479.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1656.830 2964.800 1659.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1836.830 2964.800 1839.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2016.830 2964.800 2019.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2196.830 2964.800 2199.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2376.830 2964.800 2379.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2556.830 2964.800 2559.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2736.830 2964.800 2739.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2916.830 2964.800 2919.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3096.830 2964.800 3099.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3276.830 2964.800 3279.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3456.830 2964.800 3459.930 ;
    END
    PORT
      LAYER met5 ;
        RECT 31.470 448.950 754.570 452.050 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -25.980 -20.620 -22.880 3540.300 ;
    END
    PORT
      LAYER met5 ;
        RECT -25.980 -20.620 2945.600 -17.520 ;
    END
    PORT
      LAYER met5 ;
        RECT -25.980 3537.200 2945.600 3540.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 2942.500 -20.620 2945.600 3540.300 ;
    END
    PORT
      LAYER met4 ;
        RECT 76.470 -39.820 79.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 256.470 -39.820 259.570 167.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 256.470 1006.000 259.570 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 256.470 3352.380 259.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 436.470 -39.820 439.570 167.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 436.470 1006.000 439.570 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 436.470 3352.380 439.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 616.470 -39.820 619.570 167.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 616.470 1006.000 619.570 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 616.470 3352.380 619.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 796.470 -39.820 799.570 567.420 ;
    END
    PORT
      LAYER met4 ;
        RECT 796.470 1006.000 799.570 1464.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 796.470 2157.140 799.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 976.470 -39.820 979.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1156.470 -39.820 1159.570 990.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1156.470 1247.250 1159.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1336.470 -39.820 1339.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1516.470 -39.820 1519.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1696.470 -39.820 1699.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1696.470 2742.900 1699.570 3018.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1696.470 3365.040 1699.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 1876.470 -39.820 1879.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1876.470 2742.900 1879.570 3018.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 1876.470 3365.040 1879.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2056.470 -39.820 2059.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2056.470 2742.900 2059.570 3018.940 ;
    END
    PORT
      LAYER met4 ;
        RECT 2056.470 3365.040 2059.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2236.470 -39.820 2239.570 786.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2236.470 1224.580 2239.570 2050.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 2236.470 2742.900 2239.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2416.470 -39.820 2419.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2416.470 613.620 2419.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2596.470 -39.820 2599.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2596.470 613.620 2599.570 3559.500 ;
    END
    PORT
      LAYER met4 ;
        RECT 2776.470 -39.820 2779.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2776.470 613.620 2779.570 3559.500 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 81.830 2964.800 84.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 261.830 2964.800 264.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 441.830 2964.800 444.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 621.830 2964.800 624.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 801.830 2964.800 804.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 981.830 2964.800 984.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1161.830 2964.800 1164.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1341.830 2964.800 1344.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1521.830 2964.800 1524.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1701.830 2964.800 1704.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 1881.830 2964.800 1884.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2061.830 2964.800 2064.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2241.830 2964.800 2244.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2421.830 2964.800 2424.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2601.830 2964.800 2604.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2781.830 2964.800 2784.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 2961.830 2964.800 2964.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3141.830 2964.800 3144.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3321.830 2964.800 3324.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -45.180 3501.830 2964.800 3504.930 ;
    END
  END vssd2
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.850 -4.800 99.410 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.370 -4.800 104.930 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.890 -4.800 110.450 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.970 -4.800 132.530 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.650 -4.800 320.210 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 336.210 -4.800 336.770 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.770 -4.800 353.330 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 369.330 -4.800 369.890 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.890 -4.800 386.450 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.450 -4.800 403.010 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 419.010 -4.800 419.570 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.570 -4.800 436.130 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 452.130 -4.800 452.690 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.690 -4.800 469.250 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.050 -4.800 154.610 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.250 -4.800 485.810 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.810 -4.800 502.370 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.370 -4.800 518.930 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.930 -4.800 535.490 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.490 -4.800 552.050 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 568.050 -4.800 568.610 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.610 -4.800 585.170 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 601.170 -4.800 601.730 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.730 -4.800 618.290 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.290 -4.800 634.850 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 176.130 -4.800 176.690 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.410 -4.800 667.970 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.210 -4.800 198.770 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 220.290 -4.800 220.850 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.850 -4.800 237.410 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.410 -4.800 253.970 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.970 -4.800 270.530 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.530 -4.800 287.090 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.090 -4.800 303.650 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.410 -4.800 115.970 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.490 -4.800 138.050 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.170 -4.800 325.730 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.730 -4.800 342.290 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 358.290 -4.800 358.850 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.850 -4.800 375.410 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 391.410 -4.800 391.970 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.970 -4.800 408.530 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.530 -4.800 425.090 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 441.090 -4.800 441.650 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.650 -4.800 458.210 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 474.210 -4.800 474.770 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.570 -4.800 160.130 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.770 -4.800 491.330 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 507.330 -4.800 507.890 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.890 -4.800 524.450 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.450 -4.800 541.010 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.010 -4.800 557.570 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.570 -4.800 574.130 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.130 -4.800 590.690 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.690 -4.800 607.250 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.250 -4.800 623.810 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.810 -4.800 640.370 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.650 -4.800 182.210 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 656.370 -4.800 656.930 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.930 -4.800 673.490 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.730 -4.800 204.290 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.810 -4.800 226.370 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.370 -4.800 242.930 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.930 -4.800 259.490 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.490 -4.800 276.050 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.050 -4.800 292.610 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.610 -4.800 309.170 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.010 -4.800 143.570 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.690 -4.800 331.250 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.250 -4.800 347.810 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.810 -4.800 364.370 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.370 -4.800 380.930 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.930 -4.800 397.490 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.490 -4.800 414.050 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 430.050 -4.800 430.610 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.610 -4.800 447.170 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.170 -4.800 463.730 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.730 -4.800 480.290 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.090 -4.800 165.650 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 496.290 -4.800 496.850 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.850 -4.800 513.410 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 529.410 -4.800 529.970 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.970 -4.800 546.530 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.530 -4.800 563.090 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.090 -4.800 579.650 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.650 -4.800 596.210 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.210 -4.800 612.770 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.770 -4.800 629.330 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.330 -4.800 645.890 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 187.170 -4.800 187.730 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.890 -4.800 662.450 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.450 -4.800 679.010 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.250 -4.800 209.810 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.330 -4.800 231.890 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.890 -4.800 248.450 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.450 -4.800 265.010 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.010 -4.800 281.570 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.570 -4.800 298.130 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.130 -4.800 314.690 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.530 -4.800 149.090 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.610 -4.800 171.170 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.690 -4.800 193.250 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.770 -4.800 215.330 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.930 -4.800 121.490 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.450 -4.800 127.010 2.400 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2914.100 3508.885 ;
      LAYER met1 ;
        RECT 5.520 1.740 2914.570 3515.220 ;
      LAYER met2 ;
        RECT 6.990 3517.320 42.450 3518.050 ;
        RECT 43.570 3517.320 123.410 3518.050 ;
        RECT 124.530 3517.320 204.370 3518.050 ;
        RECT 205.490 3517.320 285.330 3518.050 ;
        RECT 286.450 3517.320 366.290 3518.050 ;
        RECT 367.410 3517.320 447.250 3518.050 ;
        RECT 448.370 3517.320 528.210 3518.050 ;
        RECT 529.330 3517.320 609.170 3518.050 ;
        RECT 610.290 3517.320 690.130 3518.050 ;
        RECT 691.250 3517.320 771.090 3518.050 ;
        RECT 772.210 3517.320 852.050 3518.050 ;
        RECT 853.170 3517.320 933.010 3518.050 ;
        RECT 934.130 3517.320 1013.970 3518.050 ;
        RECT 1015.090 3517.320 1094.930 3518.050 ;
        RECT 1096.050 3517.320 1175.890 3518.050 ;
        RECT 1177.010 3517.320 1256.850 3518.050 ;
        RECT 1257.970 3517.320 1337.810 3518.050 ;
        RECT 1338.930 3517.320 1418.770 3518.050 ;
        RECT 1419.890 3517.320 1499.730 3518.050 ;
        RECT 1500.850 3517.320 1580.690 3518.050 ;
        RECT 1581.810 3517.320 1661.650 3518.050 ;
        RECT 1662.770 3517.320 1742.610 3518.050 ;
        RECT 1743.730 3517.320 1823.570 3518.050 ;
        RECT 1824.690 3517.320 1904.530 3518.050 ;
        RECT 1905.650 3517.320 1985.490 3518.050 ;
        RECT 1986.610 3517.320 2066.450 3518.050 ;
        RECT 2067.570 3517.320 2147.410 3518.050 ;
        RECT 2148.530 3517.320 2228.370 3518.050 ;
        RECT 2229.490 3517.320 2309.330 3518.050 ;
        RECT 2310.450 3517.320 2390.290 3518.050 ;
        RECT 2391.410 3517.320 2471.250 3518.050 ;
        RECT 2472.370 3517.320 2552.210 3518.050 ;
        RECT 2553.330 3517.320 2633.170 3518.050 ;
        RECT 2634.290 3517.320 2714.130 3518.050 ;
        RECT 2715.250 3517.320 2795.090 3518.050 ;
        RECT 2796.210 3517.320 2876.050 3518.050 ;
        RECT 2877.170 3517.320 2914.430 3518.050 ;
        RECT 6.990 2.680 2914.430 3517.320 ;
        RECT 6.990 1.630 98.570 2.680 ;
        RECT 99.690 1.630 104.090 2.680 ;
        RECT 105.210 1.630 109.610 2.680 ;
        RECT 110.730 1.630 115.130 2.680 ;
        RECT 116.250 1.630 120.650 2.680 ;
        RECT 121.770 1.630 126.170 2.680 ;
        RECT 127.290 1.630 131.690 2.680 ;
        RECT 132.810 1.630 137.210 2.680 ;
        RECT 138.330 1.630 142.730 2.680 ;
        RECT 143.850 1.630 148.250 2.680 ;
        RECT 149.370 1.630 153.770 2.680 ;
        RECT 154.890 1.630 159.290 2.680 ;
        RECT 160.410 1.630 164.810 2.680 ;
        RECT 165.930 1.630 170.330 2.680 ;
        RECT 171.450 1.630 175.850 2.680 ;
        RECT 176.970 1.630 181.370 2.680 ;
        RECT 182.490 1.630 186.890 2.680 ;
        RECT 188.010 1.630 192.410 2.680 ;
        RECT 193.530 1.630 197.930 2.680 ;
        RECT 199.050 1.630 203.450 2.680 ;
        RECT 204.570 1.630 208.970 2.680 ;
        RECT 210.090 1.630 214.490 2.680 ;
        RECT 215.610 1.630 220.010 2.680 ;
        RECT 221.130 1.630 225.530 2.680 ;
        RECT 226.650 1.630 231.050 2.680 ;
        RECT 232.170 1.630 236.570 2.680 ;
        RECT 237.690 1.630 242.090 2.680 ;
        RECT 243.210 1.630 247.610 2.680 ;
        RECT 248.730 1.630 253.130 2.680 ;
        RECT 254.250 1.630 258.650 2.680 ;
        RECT 259.770 1.630 264.170 2.680 ;
        RECT 265.290 1.630 269.690 2.680 ;
        RECT 270.810 1.630 275.210 2.680 ;
        RECT 276.330 1.630 280.730 2.680 ;
        RECT 281.850 1.630 286.250 2.680 ;
        RECT 287.370 1.630 291.770 2.680 ;
        RECT 292.890 1.630 297.290 2.680 ;
        RECT 298.410 1.630 302.810 2.680 ;
        RECT 303.930 1.630 308.330 2.680 ;
        RECT 309.450 1.630 313.850 2.680 ;
        RECT 314.970 1.630 319.370 2.680 ;
        RECT 320.490 1.630 324.890 2.680 ;
        RECT 326.010 1.630 330.410 2.680 ;
        RECT 331.530 1.630 335.930 2.680 ;
        RECT 337.050 1.630 341.450 2.680 ;
        RECT 342.570 1.630 346.970 2.680 ;
        RECT 348.090 1.630 352.490 2.680 ;
        RECT 353.610 1.630 358.010 2.680 ;
        RECT 359.130 1.630 363.530 2.680 ;
        RECT 364.650 1.630 369.050 2.680 ;
        RECT 370.170 1.630 374.570 2.680 ;
        RECT 375.690 1.630 380.090 2.680 ;
        RECT 381.210 1.630 385.610 2.680 ;
        RECT 386.730 1.630 391.130 2.680 ;
        RECT 392.250 1.630 396.650 2.680 ;
        RECT 397.770 1.630 402.170 2.680 ;
        RECT 403.290 1.630 407.690 2.680 ;
        RECT 408.810 1.630 413.210 2.680 ;
        RECT 414.330 1.630 418.730 2.680 ;
        RECT 419.850 1.630 424.250 2.680 ;
        RECT 425.370 1.630 429.770 2.680 ;
        RECT 430.890 1.630 435.290 2.680 ;
        RECT 436.410 1.630 440.810 2.680 ;
        RECT 441.930 1.630 446.330 2.680 ;
        RECT 447.450 1.630 451.850 2.680 ;
        RECT 452.970 1.630 457.370 2.680 ;
        RECT 458.490 1.630 462.890 2.680 ;
        RECT 464.010 1.630 468.410 2.680 ;
        RECT 469.530 1.630 473.930 2.680 ;
        RECT 475.050 1.630 479.450 2.680 ;
        RECT 480.570 1.630 484.970 2.680 ;
        RECT 486.090 1.630 490.490 2.680 ;
        RECT 491.610 1.630 496.010 2.680 ;
        RECT 497.130 1.630 501.530 2.680 ;
        RECT 502.650 1.630 507.050 2.680 ;
        RECT 508.170 1.630 512.570 2.680 ;
        RECT 513.690 1.630 518.090 2.680 ;
        RECT 519.210 1.630 523.610 2.680 ;
        RECT 524.730 1.630 529.130 2.680 ;
        RECT 530.250 1.630 534.650 2.680 ;
        RECT 535.770 1.630 540.170 2.680 ;
        RECT 541.290 1.630 545.690 2.680 ;
        RECT 546.810 1.630 551.210 2.680 ;
        RECT 552.330 1.630 556.730 2.680 ;
        RECT 557.850 1.630 562.250 2.680 ;
        RECT 563.370 1.630 567.770 2.680 ;
        RECT 568.890 1.630 573.290 2.680 ;
        RECT 574.410 1.630 578.810 2.680 ;
        RECT 579.930 1.630 584.330 2.680 ;
        RECT 585.450 1.630 589.850 2.680 ;
        RECT 590.970 1.630 595.370 2.680 ;
        RECT 596.490 1.630 600.890 2.680 ;
        RECT 602.010 1.630 606.410 2.680 ;
        RECT 607.530 1.630 611.930 2.680 ;
        RECT 613.050 1.630 617.450 2.680 ;
        RECT 618.570 1.630 622.970 2.680 ;
        RECT 624.090 1.630 628.490 2.680 ;
        RECT 629.610 1.630 634.010 2.680 ;
        RECT 635.130 1.630 639.530 2.680 ;
        RECT 640.650 1.630 645.050 2.680 ;
        RECT 646.170 1.630 650.570 2.680 ;
        RECT 651.690 1.630 656.090 2.680 ;
        RECT 657.210 1.630 661.610 2.680 ;
        RECT 662.730 1.630 667.130 2.680 ;
        RECT 668.250 1.630 672.650 2.680 ;
        RECT 673.770 1.630 678.170 2.680 ;
        RECT 679.290 1.630 683.690 2.680 ;
        RECT 684.810 1.630 689.210 2.680 ;
        RECT 690.330 1.630 694.730 2.680 ;
        RECT 695.850 1.630 700.250 2.680 ;
        RECT 701.370 1.630 705.770 2.680 ;
        RECT 706.890 1.630 711.290 2.680 ;
        RECT 712.410 1.630 716.810 2.680 ;
        RECT 717.930 1.630 722.330 2.680 ;
        RECT 723.450 1.630 727.850 2.680 ;
        RECT 728.970 1.630 733.370 2.680 ;
        RECT 734.490 1.630 738.890 2.680 ;
        RECT 740.010 1.630 744.410 2.680 ;
        RECT 745.530 1.630 749.930 2.680 ;
        RECT 751.050 1.630 755.450 2.680 ;
        RECT 756.570 1.630 760.970 2.680 ;
        RECT 762.090 1.630 766.490 2.680 ;
        RECT 767.610 1.630 772.010 2.680 ;
        RECT 773.130 1.630 777.530 2.680 ;
        RECT 778.650 1.630 783.050 2.680 ;
        RECT 784.170 1.630 788.570 2.680 ;
        RECT 789.690 1.630 794.090 2.680 ;
        RECT 795.210 1.630 799.610 2.680 ;
        RECT 800.730 1.630 805.130 2.680 ;
        RECT 806.250 1.630 810.650 2.680 ;
        RECT 811.770 1.630 816.170 2.680 ;
        RECT 817.290 1.630 821.690 2.680 ;
        RECT 822.810 1.630 827.210 2.680 ;
        RECT 828.330 1.630 832.730 2.680 ;
        RECT 833.850 1.630 838.250 2.680 ;
        RECT 839.370 1.630 843.770 2.680 ;
        RECT 844.890 1.630 849.290 2.680 ;
        RECT 850.410 1.630 854.810 2.680 ;
        RECT 855.930 1.630 860.330 2.680 ;
        RECT 861.450 1.630 865.850 2.680 ;
        RECT 866.970 1.630 871.370 2.680 ;
        RECT 872.490 1.630 876.890 2.680 ;
        RECT 878.010 1.630 882.410 2.680 ;
        RECT 883.530 1.630 887.930 2.680 ;
        RECT 889.050 1.630 893.450 2.680 ;
        RECT 894.570 1.630 898.970 2.680 ;
        RECT 900.090 1.630 904.490 2.680 ;
        RECT 905.610 1.630 910.010 2.680 ;
        RECT 911.130 1.630 915.530 2.680 ;
        RECT 916.650 1.630 921.050 2.680 ;
        RECT 922.170 1.630 926.570 2.680 ;
        RECT 927.690 1.630 932.090 2.680 ;
        RECT 933.210 1.630 937.610 2.680 ;
        RECT 938.730 1.630 943.130 2.680 ;
        RECT 944.250 1.630 948.650 2.680 ;
        RECT 949.770 1.630 954.170 2.680 ;
        RECT 955.290 1.630 959.690 2.680 ;
        RECT 960.810 1.630 965.210 2.680 ;
        RECT 966.330 1.630 970.730 2.680 ;
        RECT 971.850 1.630 976.250 2.680 ;
        RECT 977.370 1.630 981.770 2.680 ;
        RECT 982.890 1.630 987.290 2.680 ;
        RECT 988.410 1.630 992.810 2.680 ;
        RECT 993.930 1.630 998.330 2.680 ;
        RECT 999.450 1.630 1003.850 2.680 ;
        RECT 1004.970 1.630 1009.370 2.680 ;
        RECT 1010.490 1.630 1014.890 2.680 ;
        RECT 1016.010 1.630 1020.410 2.680 ;
        RECT 1021.530 1.630 1025.930 2.680 ;
        RECT 1027.050 1.630 1031.450 2.680 ;
        RECT 1032.570 1.630 1036.970 2.680 ;
        RECT 1038.090 1.630 1042.490 2.680 ;
        RECT 1043.610 1.630 1048.010 2.680 ;
        RECT 1049.130 1.630 1053.530 2.680 ;
        RECT 1054.650 1.630 1059.050 2.680 ;
        RECT 1060.170 1.630 1064.570 2.680 ;
        RECT 1065.690 1.630 1070.090 2.680 ;
        RECT 1071.210 1.630 1075.610 2.680 ;
        RECT 1076.730 1.630 1081.130 2.680 ;
        RECT 1082.250 1.630 1086.650 2.680 ;
        RECT 1087.770 1.630 1092.170 2.680 ;
        RECT 1093.290 1.630 1097.690 2.680 ;
        RECT 1098.810 1.630 1103.210 2.680 ;
        RECT 1104.330 1.630 1108.730 2.680 ;
        RECT 1109.850 1.630 1114.250 2.680 ;
        RECT 1115.370 1.630 1119.770 2.680 ;
        RECT 1120.890 1.630 1125.290 2.680 ;
        RECT 1126.410 1.630 1130.810 2.680 ;
        RECT 1131.930 1.630 1136.330 2.680 ;
        RECT 1137.450 1.630 1141.850 2.680 ;
        RECT 1142.970 1.630 1147.370 2.680 ;
        RECT 1148.490 1.630 1152.890 2.680 ;
        RECT 1154.010 1.630 1158.410 2.680 ;
        RECT 1159.530 1.630 1163.930 2.680 ;
        RECT 1165.050 1.630 1169.450 2.680 ;
        RECT 1170.570 1.630 1174.970 2.680 ;
        RECT 1176.090 1.630 1180.490 2.680 ;
        RECT 1181.610 1.630 1186.010 2.680 ;
        RECT 1187.130 1.630 1191.530 2.680 ;
        RECT 1192.650 1.630 1197.050 2.680 ;
        RECT 1198.170 1.630 1202.570 2.680 ;
        RECT 1203.690 1.630 1208.090 2.680 ;
        RECT 1209.210 1.630 1213.610 2.680 ;
        RECT 1214.730 1.630 1219.130 2.680 ;
        RECT 1220.250 1.630 1224.650 2.680 ;
        RECT 1225.770 1.630 1230.170 2.680 ;
        RECT 1231.290 1.630 1235.690 2.680 ;
        RECT 1236.810 1.630 1241.210 2.680 ;
        RECT 1242.330 1.630 1246.730 2.680 ;
        RECT 1247.850 1.630 1252.250 2.680 ;
        RECT 1253.370 1.630 1257.770 2.680 ;
        RECT 1258.890 1.630 1263.290 2.680 ;
        RECT 1264.410 1.630 1268.810 2.680 ;
        RECT 1269.930 1.630 1274.330 2.680 ;
        RECT 1275.450 1.630 1279.850 2.680 ;
        RECT 1280.970 1.630 1285.370 2.680 ;
        RECT 1286.490 1.630 1290.890 2.680 ;
        RECT 1292.010 1.630 1296.410 2.680 ;
        RECT 1297.530 1.630 1301.930 2.680 ;
        RECT 1303.050 1.630 1307.450 2.680 ;
        RECT 1308.570 1.630 1312.970 2.680 ;
        RECT 1314.090 1.630 1318.490 2.680 ;
        RECT 1319.610 1.630 1324.010 2.680 ;
        RECT 1325.130 1.630 1329.530 2.680 ;
        RECT 1330.650 1.630 1335.050 2.680 ;
        RECT 1336.170 1.630 1340.570 2.680 ;
        RECT 1341.690 1.630 1346.090 2.680 ;
        RECT 1347.210 1.630 1351.610 2.680 ;
        RECT 1352.730 1.630 1357.130 2.680 ;
        RECT 1358.250 1.630 1362.650 2.680 ;
        RECT 1363.770 1.630 1368.170 2.680 ;
        RECT 1369.290 1.630 1373.690 2.680 ;
        RECT 1374.810 1.630 1379.210 2.680 ;
        RECT 1380.330 1.630 1384.730 2.680 ;
        RECT 1385.850 1.630 1390.250 2.680 ;
        RECT 1391.370 1.630 1395.770 2.680 ;
        RECT 1396.890 1.630 1401.290 2.680 ;
        RECT 1402.410 1.630 1406.810 2.680 ;
        RECT 1407.930 1.630 1412.330 2.680 ;
        RECT 1413.450 1.630 1417.850 2.680 ;
        RECT 1418.970 1.630 1423.370 2.680 ;
        RECT 1424.490 1.630 1428.890 2.680 ;
        RECT 1430.010 1.630 1434.410 2.680 ;
        RECT 1435.530 1.630 1439.930 2.680 ;
        RECT 1441.050 1.630 1445.450 2.680 ;
        RECT 1446.570 1.630 1450.970 2.680 ;
        RECT 1452.090 1.630 1456.490 2.680 ;
        RECT 1457.610 1.630 1462.010 2.680 ;
        RECT 1463.130 1.630 1467.530 2.680 ;
        RECT 1468.650 1.630 1473.050 2.680 ;
        RECT 1474.170 1.630 1478.570 2.680 ;
        RECT 1479.690 1.630 1484.090 2.680 ;
        RECT 1485.210 1.630 1489.610 2.680 ;
        RECT 1490.730 1.630 1495.130 2.680 ;
        RECT 1496.250 1.630 1500.650 2.680 ;
        RECT 1501.770 1.630 1506.170 2.680 ;
        RECT 1507.290 1.630 1511.690 2.680 ;
        RECT 1512.810 1.630 1517.210 2.680 ;
        RECT 1518.330 1.630 1522.730 2.680 ;
        RECT 1523.850 1.630 1528.250 2.680 ;
        RECT 1529.370 1.630 1533.770 2.680 ;
        RECT 1534.890 1.630 1539.290 2.680 ;
        RECT 1540.410 1.630 1544.810 2.680 ;
        RECT 1545.930 1.630 1550.330 2.680 ;
        RECT 1551.450 1.630 1555.850 2.680 ;
        RECT 1556.970 1.630 1561.370 2.680 ;
        RECT 1562.490 1.630 1566.890 2.680 ;
        RECT 1568.010 1.630 1572.410 2.680 ;
        RECT 1573.530 1.630 1577.930 2.680 ;
        RECT 1579.050 1.630 1583.450 2.680 ;
        RECT 1584.570 1.630 1588.970 2.680 ;
        RECT 1590.090 1.630 1594.490 2.680 ;
        RECT 1595.610 1.630 1600.010 2.680 ;
        RECT 1601.130 1.630 1605.530 2.680 ;
        RECT 1606.650 1.630 1611.050 2.680 ;
        RECT 1612.170 1.630 1616.570 2.680 ;
        RECT 1617.690 1.630 1622.090 2.680 ;
        RECT 1623.210 1.630 1627.610 2.680 ;
        RECT 1628.730 1.630 1633.130 2.680 ;
        RECT 1634.250 1.630 1638.650 2.680 ;
        RECT 1639.770 1.630 1644.170 2.680 ;
        RECT 1645.290 1.630 1649.690 2.680 ;
        RECT 1650.810 1.630 1655.210 2.680 ;
        RECT 1656.330 1.630 1660.730 2.680 ;
        RECT 1661.850 1.630 1666.250 2.680 ;
        RECT 1667.370 1.630 1671.770 2.680 ;
        RECT 1672.890 1.630 1677.290 2.680 ;
        RECT 1678.410 1.630 1682.810 2.680 ;
        RECT 1683.930 1.630 1688.330 2.680 ;
        RECT 1689.450 1.630 1693.850 2.680 ;
        RECT 1694.970 1.630 1699.370 2.680 ;
        RECT 1700.490 1.630 1704.890 2.680 ;
        RECT 1706.010 1.630 1710.410 2.680 ;
        RECT 1711.530 1.630 1715.930 2.680 ;
        RECT 1717.050 1.630 1721.450 2.680 ;
        RECT 1722.570 1.630 1726.970 2.680 ;
        RECT 1728.090 1.630 1732.490 2.680 ;
        RECT 1733.610 1.630 1738.010 2.680 ;
        RECT 1739.130 1.630 1743.530 2.680 ;
        RECT 1744.650 1.630 1749.050 2.680 ;
        RECT 1750.170 1.630 1754.570 2.680 ;
        RECT 1755.690 1.630 1760.090 2.680 ;
        RECT 1761.210 1.630 1765.610 2.680 ;
        RECT 1766.730 1.630 1771.130 2.680 ;
        RECT 1772.250 1.630 1776.650 2.680 ;
        RECT 1777.770 1.630 1782.170 2.680 ;
        RECT 1783.290 1.630 1787.690 2.680 ;
        RECT 1788.810 1.630 1793.210 2.680 ;
        RECT 1794.330 1.630 1798.730 2.680 ;
        RECT 1799.850 1.630 1804.250 2.680 ;
        RECT 1805.370 1.630 1809.770 2.680 ;
        RECT 1810.890 1.630 1815.290 2.680 ;
        RECT 1816.410 1.630 1820.810 2.680 ;
        RECT 1821.930 1.630 1826.330 2.680 ;
        RECT 1827.450 1.630 1831.850 2.680 ;
        RECT 1832.970 1.630 1837.370 2.680 ;
        RECT 1838.490 1.630 1842.890 2.680 ;
        RECT 1844.010 1.630 1848.410 2.680 ;
        RECT 1849.530 1.630 1853.930 2.680 ;
        RECT 1855.050 1.630 1859.450 2.680 ;
        RECT 1860.570 1.630 1864.970 2.680 ;
        RECT 1866.090 1.630 1870.490 2.680 ;
        RECT 1871.610 1.630 1876.010 2.680 ;
        RECT 1877.130 1.630 1881.530 2.680 ;
        RECT 1882.650 1.630 1887.050 2.680 ;
        RECT 1888.170 1.630 1892.570 2.680 ;
        RECT 1893.690 1.630 1898.090 2.680 ;
        RECT 1899.210 1.630 1903.610 2.680 ;
        RECT 1904.730 1.630 1909.130 2.680 ;
        RECT 1910.250 1.630 1914.650 2.680 ;
        RECT 1915.770 1.630 1920.170 2.680 ;
        RECT 1921.290 1.630 1925.690 2.680 ;
        RECT 1926.810 1.630 1931.210 2.680 ;
        RECT 1932.330 1.630 1936.730 2.680 ;
        RECT 1937.850 1.630 1942.250 2.680 ;
        RECT 1943.370 1.630 1947.770 2.680 ;
        RECT 1948.890 1.630 1953.290 2.680 ;
        RECT 1954.410 1.630 1958.810 2.680 ;
        RECT 1959.930 1.630 1964.330 2.680 ;
        RECT 1965.450 1.630 1969.850 2.680 ;
        RECT 1970.970 1.630 1975.370 2.680 ;
        RECT 1976.490 1.630 1980.890 2.680 ;
        RECT 1982.010 1.630 1986.410 2.680 ;
        RECT 1987.530 1.630 1991.930 2.680 ;
        RECT 1993.050 1.630 1997.450 2.680 ;
        RECT 1998.570 1.630 2002.970 2.680 ;
        RECT 2004.090 1.630 2008.490 2.680 ;
        RECT 2009.610 1.630 2014.010 2.680 ;
        RECT 2015.130 1.630 2019.530 2.680 ;
        RECT 2020.650 1.630 2025.050 2.680 ;
        RECT 2026.170 1.630 2030.570 2.680 ;
        RECT 2031.690 1.630 2036.090 2.680 ;
        RECT 2037.210 1.630 2041.610 2.680 ;
        RECT 2042.730 1.630 2047.130 2.680 ;
        RECT 2048.250 1.630 2052.650 2.680 ;
        RECT 2053.770 1.630 2058.170 2.680 ;
        RECT 2059.290 1.630 2063.690 2.680 ;
        RECT 2064.810 1.630 2069.210 2.680 ;
        RECT 2070.330 1.630 2074.730 2.680 ;
        RECT 2075.850 1.630 2080.250 2.680 ;
        RECT 2081.370 1.630 2085.770 2.680 ;
        RECT 2086.890 1.630 2091.290 2.680 ;
        RECT 2092.410 1.630 2096.810 2.680 ;
        RECT 2097.930 1.630 2102.330 2.680 ;
        RECT 2103.450 1.630 2107.850 2.680 ;
        RECT 2108.970 1.630 2113.370 2.680 ;
        RECT 2114.490 1.630 2118.890 2.680 ;
        RECT 2120.010 1.630 2124.410 2.680 ;
        RECT 2125.530 1.630 2129.930 2.680 ;
        RECT 2131.050 1.630 2135.450 2.680 ;
        RECT 2136.570 1.630 2140.970 2.680 ;
        RECT 2142.090 1.630 2146.490 2.680 ;
        RECT 2147.610 1.630 2152.010 2.680 ;
        RECT 2153.130 1.630 2157.530 2.680 ;
        RECT 2158.650 1.630 2163.050 2.680 ;
        RECT 2164.170 1.630 2168.570 2.680 ;
        RECT 2169.690 1.630 2174.090 2.680 ;
        RECT 2175.210 1.630 2179.610 2.680 ;
        RECT 2180.730 1.630 2185.130 2.680 ;
        RECT 2186.250 1.630 2190.650 2.680 ;
        RECT 2191.770 1.630 2196.170 2.680 ;
        RECT 2197.290 1.630 2201.690 2.680 ;
        RECT 2202.810 1.630 2207.210 2.680 ;
        RECT 2208.330 1.630 2212.730 2.680 ;
        RECT 2213.850 1.630 2218.250 2.680 ;
        RECT 2219.370 1.630 2223.770 2.680 ;
        RECT 2224.890 1.630 2229.290 2.680 ;
        RECT 2230.410 1.630 2234.810 2.680 ;
        RECT 2235.930 1.630 2240.330 2.680 ;
        RECT 2241.450 1.630 2245.850 2.680 ;
        RECT 2246.970 1.630 2251.370 2.680 ;
        RECT 2252.490 1.630 2256.890 2.680 ;
        RECT 2258.010 1.630 2262.410 2.680 ;
        RECT 2263.530 1.630 2267.930 2.680 ;
        RECT 2269.050 1.630 2273.450 2.680 ;
        RECT 2274.570 1.630 2278.970 2.680 ;
        RECT 2280.090 1.630 2284.490 2.680 ;
        RECT 2285.610 1.630 2290.010 2.680 ;
        RECT 2291.130 1.630 2295.530 2.680 ;
        RECT 2296.650 1.630 2301.050 2.680 ;
        RECT 2302.170 1.630 2306.570 2.680 ;
        RECT 2307.690 1.630 2312.090 2.680 ;
        RECT 2313.210 1.630 2317.610 2.680 ;
        RECT 2318.730 1.630 2323.130 2.680 ;
        RECT 2324.250 1.630 2328.650 2.680 ;
        RECT 2329.770 1.630 2334.170 2.680 ;
        RECT 2335.290 1.630 2339.690 2.680 ;
        RECT 2340.810 1.630 2345.210 2.680 ;
        RECT 2346.330 1.630 2350.730 2.680 ;
        RECT 2351.850 1.630 2356.250 2.680 ;
        RECT 2357.370 1.630 2361.770 2.680 ;
        RECT 2362.890 1.630 2367.290 2.680 ;
        RECT 2368.410 1.630 2372.810 2.680 ;
        RECT 2373.930 1.630 2378.330 2.680 ;
        RECT 2379.450 1.630 2383.850 2.680 ;
        RECT 2384.970 1.630 2389.370 2.680 ;
        RECT 2390.490 1.630 2394.890 2.680 ;
        RECT 2396.010 1.630 2400.410 2.680 ;
        RECT 2401.530 1.630 2405.930 2.680 ;
        RECT 2407.050 1.630 2411.450 2.680 ;
        RECT 2412.570 1.630 2416.970 2.680 ;
        RECT 2418.090 1.630 2422.490 2.680 ;
        RECT 2423.610 1.630 2428.010 2.680 ;
        RECT 2429.130 1.630 2433.530 2.680 ;
        RECT 2434.650 1.630 2439.050 2.680 ;
        RECT 2440.170 1.630 2444.570 2.680 ;
        RECT 2445.690 1.630 2450.090 2.680 ;
        RECT 2451.210 1.630 2455.610 2.680 ;
        RECT 2456.730 1.630 2461.130 2.680 ;
        RECT 2462.250 1.630 2466.650 2.680 ;
        RECT 2467.770 1.630 2472.170 2.680 ;
        RECT 2473.290 1.630 2477.690 2.680 ;
        RECT 2478.810 1.630 2483.210 2.680 ;
        RECT 2484.330 1.630 2488.730 2.680 ;
        RECT 2489.850 1.630 2494.250 2.680 ;
        RECT 2495.370 1.630 2499.770 2.680 ;
        RECT 2500.890 1.630 2505.290 2.680 ;
        RECT 2506.410 1.630 2510.810 2.680 ;
        RECT 2511.930 1.630 2516.330 2.680 ;
        RECT 2517.450 1.630 2521.850 2.680 ;
        RECT 2522.970 1.630 2527.370 2.680 ;
        RECT 2528.490 1.630 2532.890 2.680 ;
        RECT 2534.010 1.630 2538.410 2.680 ;
        RECT 2539.530 1.630 2543.930 2.680 ;
        RECT 2545.050 1.630 2549.450 2.680 ;
        RECT 2550.570 1.630 2554.970 2.680 ;
        RECT 2556.090 1.630 2560.490 2.680 ;
        RECT 2561.610 1.630 2566.010 2.680 ;
        RECT 2567.130 1.630 2571.530 2.680 ;
        RECT 2572.650 1.630 2577.050 2.680 ;
        RECT 2578.170 1.630 2582.570 2.680 ;
        RECT 2583.690 1.630 2588.090 2.680 ;
        RECT 2589.210 1.630 2593.610 2.680 ;
        RECT 2594.730 1.630 2599.130 2.680 ;
        RECT 2600.250 1.630 2604.650 2.680 ;
        RECT 2605.770 1.630 2610.170 2.680 ;
        RECT 2611.290 1.630 2615.690 2.680 ;
        RECT 2616.810 1.630 2621.210 2.680 ;
        RECT 2622.330 1.630 2626.730 2.680 ;
        RECT 2627.850 1.630 2632.250 2.680 ;
        RECT 2633.370 1.630 2637.770 2.680 ;
        RECT 2638.890 1.630 2643.290 2.680 ;
        RECT 2644.410 1.630 2648.810 2.680 ;
        RECT 2649.930 1.630 2654.330 2.680 ;
        RECT 2655.450 1.630 2659.850 2.680 ;
        RECT 2660.970 1.630 2665.370 2.680 ;
        RECT 2666.490 1.630 2670.890 2.680 ;
        RECT 2672.010 1.630 2676.410 2.680 ;
        RECT 2677.530 1.630 2681.930 2.680 ;
        RECT 2683.050 1.630 2687.450 2.680 ;
        RECT 2688.570 1.630 2692.970 2.680 ;
        RECT 2694.090 1.630 2698.490 2.680 ;
        RECT 2699.610 1.630 2704.010 2.680 ;
        RECT 2705.130 1.630 2709.530 2.680 ;
        RECT 2710.650 1.630 2715.050 2.680 ;
        RECT 2716.170 1.630 2720.570 2.680 ;
        RECT 2721.690 1.630 2726.090 2.680 ;
        RECT 2727.210 1.630 2731.610 2.680 ;
        RECT 2732.730 1.630 2737.130 2.680 ;
        RECT 2738.250 1.630 2742.650 2.680 ;
        RECT 2743.770 1.630 2748.170 2.680 ;
        RECT 2749.290 1.630 2753.690 2.680 ;
        RECT 2754.810 1.630 2759.210 2.680 ;
        RECT 2760.330 1.630 2764.730 2.680 ;
        RECT 2765.850 1.630 2770.250 2.680 ;
        RECT 2771.370 1.630 2775.770 2.680 ;
        RECT 2776.890 1.630 2781.290 2.680 ;
        RECT 2782.410 1.630 2786.810 2.680 ;
        RECT 2787.930 1.630 2792.330 2.680 ;
        RECT 2793.450 1.630 2797.850 2.680 ;
        RECT 2798.970 1.630 2803.370 2.680 ;
        RECT 2804.490 1.630 2808.890 2.680 ;
        RECT 2810.010 1.630 2814.410 2.680 ;
        RECT 2815.530 1.630 2819.930 2.680 ;
        RECT 2821.050 1.630 2914.430 2.680 ;
      LAYER met3 ;
        RECT 2.400 3475.460 2917.600 3508.965 ;
        RECT 2.400 3473.460 2917.200 3475.460 ;
        RECT 2.400 3472.740 2917.600 3473.460 ;
        RECT 2.800 3470.740 2917.600 3472.740 ;
        RECT 2.400 3409.500 2917.600 3470.740 ;
        RECT 2.400 3408.140 2917.200 3409.500 ;
        RECT 2.800 3407.500 2917.200 3408.140 ;
        RECT 2.800 3406.140 2917.600 3407.500 ;
        RECT 2.400 3343.540 2917.600 3406.140 ;
        RECT 2.800 3341.540 2917.200 3343.540 ;
        RECT 2.400 3278.940 2917.600 3341.540 ;
        RECT 2.800 3277.580 2917.600 3278.940 ;
        RECT 2.800 3276.940 2917.200 3277.580 ;
        RECT 2.400 3275.580 2917.200 3276.940 ;
        RECT 2.400 3214.340 2917.600 3275.580 ;
        RECT 2.800 3212.340 2917.600 3214.340 ;
        RECT 2.400 3211.620 2917.600 3212.340 ;
        RECT 2.400 3209.620 2917.200 3211.620 ;
        RECT 2.400 3149.740 2917.600 3209.620 ;
        RECT 2.800 3147.740 2917.600 3149.740 ;
        RECT 2.400 3145.660 2917.600 3147.740 ;
        RECT 2.400 3143.660 2917.200 3145.660 ;
        RECT 2.400 3085.140 2917.600 3143.660 ;
        RECT 2.800 3083.140 2917.600 3085.140 ;
        RECT 2.400 3079.700 2917.600 3083.140 ;
        RECT 2.400 3077.700 2917.200 3079.700 ;
        RECT 2.400 3020.540 2917.600 3077.700 ;
        RECT 2.800 3018.540 2917.600 3020.540 ;
        RECT 2.400 3013.740 2917.600 3018.540 ;
        RECT 2.400 3011.740 2917.200 3013.740 ;
        RECT 2.400 2955.940 2917.600 3011.740 ;
        RECT 2.800 2953.940 2917.600 2955.940 ;
        RECT 2.400 2947.780 2917.600 2953.940 ;
        RECT 2.400 2945.780 2917.200 2947.780 ;
        RECT 2.400 2891.340 2917.600 2945.780 ;
        RECT 2.800 2889.340 2917.600 2891.340 ;
        RECT 2.400 2881.820 2917.600 2889.340 ;
        RECT 2.400 2879.820 2917.200 2881.820 ;
        RECT 2.400 2826.740 2917.600 2879.820 ;
        RECT 2.800 2824.740 2917.600 2826.740 ;
        RECT 2.400 2815.860 2917.600 2824.740 ;
        RECT 2.400 2813.860 2917.200 2815.860 ;
        RECT 2.400 2762.140 2917.600 2813.860 ;
        RECT 2.800 2760.140 2917.600 2762.140 ;
        RECT 2.400 2749.900 2917.600 2760.140 ;
        RECT 2.400 2747.900 2917.200 2749.900 ;
        RECT 2.400 2697.540 2917.600 2747.900 ;
        RECT 2.800 2695.540 2917.600 2697.540 ;
        RECT 2.400 2683.940 2917.600 2695.540 ;
        RECT 2.400 2681.940 2917.200 2683.940 ;
        RECT 2.400 2632.940 2917.600 2681.940 ;
        RECT 2.800 2630.940 2917.600 2632.940 ;
        RECT 2.400 2617.980 2917.600 2630.940 ;
        RECT 2.400 2615.980 2917.200 2617.980 ;
        RECT 2.400 2568.340 2917.600 2615.980 ;
        RECT 2.800 2566.340 2917.600 2568.340 ;
        RECT 2.400 2552.020 2917.600 2566.340 ;
        RECT 2.400 2550.020 2917.200 2552.020 ;
        RECT 2.400 2503.740 2917.600 2550.020 ;
        RECT 2.800 2501.740 2917.600 2503.740 ;
        RECT 2.400 2486.060 2917.600 2501.740 ;
        RECT 2.400 2484.060 2917.200 2486.060 ;
        RECT 2.400 2439.140 2917.600 2484.060 ;
        RECT 2.800 2437.140 2917.600 2439.140 ;
        RECT 2.400 2420.100 2917.600 2437.140 ;
        RECT 2.400 2418.100 2917.200 2420.100 ;
        RECT 2.400 2374.540 2917.600 2418.100 ;
        RECT 2.800 2372.540 2917.600 2374.540 ;
        RECT 2.400 2354.140 2917.600 2372.540 ;
        RECT 2.400 2352.140 2917.200 2354.140 ;
        RECT 2.400 2309.940 2917.600 2352.140 ;
        RECT 2.800 2307.940 2917.600 2309.940 ;
        RECT 2.400 2288.180 2917.600 2307.940 ;
        RECT 2.400 2286.180 2917.200 2288.180 ;
        RECT 2.400 2245.340 2917.600 2286.180 ;
        RECT 2.800 2243.340 2917.600 2245.340 ;
        RECT 2.400 2222.220 2917.600 2243.340 ;
        RECT 2.400 2220.220 2917.200 2222.220 ;
        RECT 2.400 2180.740 2917.600 2220.220 ;
        RECT 2.800 2178.740 2917.600 2180.740 ;
        RECT 2.400 2156.260 2917.600 2178.740 ;
        RECT 2.400 2154.260 2917.200 2156.260 ;
        RECT 2.400 2116.140 2917.600 2154.260 ;
        RECT 2.800 2114.140 2917.600 2116.140 ;
        RECT 2.400 2090.300 2917.600 2114.140 ;
        RECT 2.400 2088.300 2917.200 2090.300 ;
        RECT 2.400 2051.540 2917.600 2088.300 ;
        RECT 2.800 2049.540 2917.600 2051.540 ;
        RECT 2.400 2024.340 2917.600 2049.540 ;
        RECT 2.400 2022.340 2917.200 2024.340 ;
        RECT 2.400 1986.940 2917.600 2022.340 ;
        RECT 2.800 1984.940 2917.600 1986.940 ;
        RECT 2.400 1958.380 2917.600 1984.940 ;
        RECT 2.400 1956.380 2917.200 1958.380 ;
        RECT 2.400 1922.340 2917.600 1956.380 ;
        RECT 2.800 1920.340 2917.600 1922.340 ;
        RECT 2.400 1892.420 2917.600 1920.340 ;
        RECT 2.400 1890.420 2917.200 1892.420 ;
        RECT 2.400 1857.740 2917.600 1890.420 ;
        RECT 2.800 1855.740 2917.600 1857.740 ;
        RECT 2.400 1826.460 2917.600 1855.740 ;
        RECT 2.400 1824.460 2917.200 1826.460 ;
        RECT 2.400 1793.140 2917.600 1824.460 ;
        RECT 2.800 1791.140 2917.600 1793.140 ;
        RECT 2.400 1760.500 2917.600 1791.140 ;
        RECT 2.400 1758.500 2917.200 1760.500 ;
        RECT 2.400 1728.540 2917.600 1758.500 ;
        RECT 2.800 1726.540 2917.600 1728.540 ;
        RECT 2.400 1694.540 2917.600 1726.540 ;
        RECT 2.400 1692.540 2917.200 1694.540 ;
        RECT 2.400 1663.940 2917.600 1692.540 ;
        RECT 2.800 1661.940 2917.600 1663.940 ;
        RECT 2.400 1628.580 2917.600 1661.940 ;
        RECT 2.400 1626.580 2917.200 1628.580 ;
        RECT 2.400 1599.340 2917.600 1626.580 ;
        RECT 2.800 1597.340 2917.600 1599.340 ;
        RECT 2.400 1562.620 2917.600 1597.340 ;
        RECT 2.400 1560.620 2917.200 1562.620 ;
        RECT 2.400 1534.740 2917.600 1560.620 ;
        RECT 2.800 1532.740 2917.600 1534.740 ;
        RECT 2.400 1496.660 2917.600 1532.740 ;
        RECT 2.400 1494.660 2917.200 1496.660 ;
        RECT 2.400 1470.140 2917.600 1494.660 ;
        RECT 2.800 1468.140 2917.600 1470.140 ;
        RECT 2.400 1430.700 2917.600 1468.140 ;
        RECT 2.400 1428.700 2917.200 1430.700 ;
        RECT 2.400 1405.540 2917.600 1428.700 ;
        RECT 2.800 1403.540 2917.600 1405.540 ;
        RECT 2.400 1364.740 2917.600 1403.540 ;
        RECT 2.400 1362.740 2917.200 1364.740 ;
        RECT 2.400 1340.940 2917.600 1362.740 ;
        RECT 2.800 1338.940 2917.600 1340.940 ;
        RECT 2.400 1298.780 2917.600 1338.940 ;
        RECT 2.400 1296.780 2917.200 1298.780 ;
        RECT 2.400 1276.340 2917.600 1296.780 ;
        RECT 2.800 1274.340 2917.600 1276.340 ;
        RECT 2.400 1232.820 2917.600 1274.340 ;
        RECT 2.400 1230.820 2917.200 1232.820 ;
        RECT 2.400 1211.740 2917.600 1230.820 ;
        RECT 2.800 1209.740 2917.600 1211.740 ;
        RECT 2.400 1166.860 2917.600 1209.740 ;
        RECT 2.400 1164.860 2917.200 1166.860 ;
        RECT 2.400 1147.140 2917.600 1164.860 ;
        RECT 2.800 1145.140 2917.600 1147.140 ;
        RECT 2.400 1100.900 2917.600 1145.140 ;
        RECT 2.400 1098.900 2917.200 1100.900 ;
        RECT 2.400 1082.540 2917.600 1098.900 ;
        RECT 2.800 1080.540 2917.600 1082.540 ;
        RECT 2.400 1034.940 2917.600 1080.540 ;
        RECT 2.400 1032.940 2917.200 1034.940 ;
        RECT 2.400 1017.940 2917.600 1032.940 ;
        RECT 2.800 1015.940 2917.600 1017.940 ;
        RECT 2.400 968.980 2917.600 1015.940 ;
        RECT 2.400 966.980 2917.200 968.980 ;
        RECT 2.400 953.340 2917.600 966.980 ;
        RECT 2.800 951.340 2917.600 953.340 ;
        RECT 2.400 903.020 2917.600 951.340 ;
        RECT 2.400 901.020 2917.200 903.020 ;
        RECT 2.400 888.740 2917.600 901.020 ;
        RECT 2.800 886.740 2917.600 888.740 ;
        RECT 2.400 837.060 2917.600 886.740 ;
        RECT 2.400 835.060 2917.200 837.060 ;
        RECT 2.400 824.140 2917.600 835.060 ;
        RECT 2.800 822.140 2917.600 824.140 ;
        RECT 2.400 771.100 2917.600 822.140 ;
        RECT 2.400 769.100 2917.200 771.100 ;
        RECT 2.400 759.540 2917.600 769.100 ;
        RECT 2.800 757.540 2917.600 759.540 ;
        RECT 2.400 705.140 2917.600 757.540 ;
        RECT 2.400 703.140 2917.200 705.140 ;
        RECT 2.400 694.940 2917.600 703.140 ;
        RECT 2.800 692.940 2917.600 694.940 ;
        RECT 2.400 639.180 2917.600 692.940 ;
        RECT 2.400 637.180 2917.200 639.180 ;
        RECT 2.400 630.340 2917.600 637.180 ;
        RECT 2.800 628.340 2917.600 630.340 ;
        RECT 2.400 573.220 2917.600 628.340 ;
        RECT 2.400 571.220 2917.200 573.220 ;
        RECT 2.400 565.740 2917.600 571.220 ;
        RECT 2.800 563.740 2917.600 565.740 ;
        RECT 2.400 507.260 2917.600 563.740 ;
        RECT 2.400 505.260 2917.200 507.260 ;
        RECT 2.400 501.140 2917.600 505.260 ;
        RECT 2.800 499.140 2917.600 501.140 ;
        RECT 2.400 441.300 2917.600 499.140 ;
        RECT 2.400 439.300 2917.200 441.300 ;
        RECT 2.400 436.540 2917.600 439.300 ;
        RECT 2.800 434.540 2917.600 436.540 ;
        RECT 2.400 375.340 2917.600 434.540 ;
        RECT 2.400 373.340 2917.200 375.340 ;
        RECT 2.400 371.940 2917.600 373.340 ;
        RECT 2.800 369.940 2917.600 371.940 ;
        RECT 2.400 309.380 2917.600 369.940 ;
        RECT 2.400 307.380 2917.200 309.380 ;
        RECT 2.400 307.340 2917.600 307.380 ;
        RECT 2.800 305.340 2917.600 307.340 ;
        RECT 2.400 243.420 2917.600 305.340 ;
        RECT 2.400 242.740 2917.200 243.420 ;
        RECT 2.800 241.420 2917.200 242.740 ;
        RECT 2.800 240.740 2917.600 241.420 ;
        RECT 2.400 178.140 2917.600 240.740 ;
        RECT 2.800 177.460 2917.600 178.140 ;
        RECT 2.800 176.140 2917.200 177.460 ;
        RECT 2.400 175.460 2917.200 176.140 ;
        RECT 2.400 113.540 2917.600 175.460 ;
        RECT 2.800 111.540 2917.600 113.540 ;
        RECT 2.400 111.500 2917.600 111.540 ;
        RECT 2.400 109.500 2917.200 111.500 ;
        RECT 2.400 48.940 2917.600 109.500 ;
        RECT 2.800 46.940 2917.600 48.940 ;
        RECT 2.400 45.540 2917.600 46.940 ;
        RECT 2.400 43.540 2917.200 45.540 ;
        RECT 2.400 4.255 2917.600 43.540 ;
      LAYER met4 ;
        RECT 180.615 3351.980 188.570 3355.040 ;
        RECT 192.470 3351.980 211.070 3355.040 ;
        RECT 214.970 3351.980 233.570 3355.040 ;
        RECT 237.470 3351.980 256.070 3355.040 ;
        RECT 259.970 3351.980 301.070 3355.040 ;
        RECT 304.970 3351.980 323.570 3355.040 ;
        RECT 327.470 3351.980 346.070 3355.040 ;
        RECT 349.970 3351.980 368.570 3355.040 ;
        RECT 372.470 3351.980 391.070 3355.040 ;
        RECT 394.970 3351.980 413.570 3355.040 ;
        RECT 417.470 3351.980 436.070 3355.040 ;
        RECT 439.970 3351.980 481.070 3355.040 ;
        RECT 484.970 3351.980 503.570 3355.040 ;
        RECT 507.470 3351.980 526.070 3355.040 ;
        RECT 529.970 3351.980 548.570 3355.040 ;
        RECT 552.470 3351.980 571.070 3355.040 ;
        RECT 574.970 3351.980 593.570 3355.040 ;
        RECT 597.470 3351.980 616.070 3355.040 ;
        RECT 619.970 3351.980 661.070 3355.040 ;
        RECT 664.970 3351.980 683.570 3355.040 ;
        RECT 180.615 2885.640 683.570 3351.980 ;
        RECT 180.615 2733.960 188.570 2885.640 ;
        RECT 192.470 2733.960 211.070 2885.640 ;
        RECT 214.970 2733.960 368.570 2885.640 ;
        RECT 372.470 2733.960 391.070 2885.640 ;
        RECT 394.970 2733.960 548.570 2885.640 ;
        RECT 552.470 2733.960 571.070 2885.640 ;
        RECT 574.970 2733.960 683.570 2885.640 ;
        RECT 687.470 2733.960 706.070 3355.040 ;
        RECT 180.615 2311.140 706.070 2733.960 ;
        RECT 180.615 2156.740 188.570 2311.140 ;
        RECT 192.470 2156.740 211.070 2311.140 ;
        RECT 214.970 2156.740 368.570 2311.140 ;
        RECT 372.470 2156.740 391.070 2311.140 ;
        RECT 394.970 2156.740 548.570 2311.140 ;
        RECT 552.470 2156.740 571.070 2311.140 ;
        RECT 574.970 2156.740 706.070 2311.140 ;
        RECT 709.970 2156.740 728.570 3355.040 ;
        RECT 732.470 2156.740 751.070 3355.040 ;
        RECT 754.970 2156.740 773.570 3355.040 ;
        RECT 777.470 2156.740 796.070 3355.040 ;
        RECT 799.970 2156.740 818.570 3355.040 ;
        RECT 822.470 2156.740 841.070 3355.040 ;
        RECT 844.970 2156.740 863.570 3355.040 ;
        RECT 867.470 2156.740 886.070 3355.040 ;
        RECT 889.970 2156.740 908.570 3355.040 ;
        RECT 912.470 2156.740 931.070 3355.040 ;
        RECT 180.615 1465.320 931.070 2156.740 ;
        RECT 180.615 1005.600 188.570 1465.320 ;
        RECT 192.470 1005.600 211.070 1465.320 ;
        RECT 214.970 1005.600 233.570 1465.320 ;
        RECT 237.470 1005.600 256.070 1465.320 ;
        RECT 259.970 1005.600 278.570 1465.320 ;
        RECT 282.470 1005.600 301.070 1465.320 ;
        RECT 304.970 1005.600 323.570 1465.320 ;
        RECT 327.470 1005.600 346.070 1465.320 ;
        RECT 349.970 1005.600 368.570 1465.320 ;
        RECT 372.470 1005.600 391.070 1465.320 ;
        RECT 394.970 1005.600 413.570 1465.320 ;
        RECT 417.470 1005.600 436.070 1465.320 ;
        RECT 439.970 1005.600 458.570 1465.320 ;
        RECT 462.470 1005.600 481.070 1465.320 ;
        RECT 484.970 1005.600 503.570 1465.320 ;
        RECT 507.470 1005.600 526.070 1465.320 ;
        RECT 529.970 1005.600 548.570 1465.320 ;
        RECT 552.470 1005.600 571.070 1465.320 ;
        RECT 574.970 1005.600 593.570 1465.320 ;
        RECT 597.470 1005.600 616.070 1465.320 ;
        RECT 619.970 1005.600 638.570 1465.320 ;
        RECT 642.470 1005.600 661.070 1465.320 ;
        RECT 664.970 1005.600 683.570 1465.320 ;
        RECT 687.470 1005.600 706.070 1465.320 ;
        RECT 709.970 1005.600 728.570 1465.320 ;
        RECT 732.470 1005.600 751.070 1465.320 ;
        RECT 754.970 1005.600 773.570 1465.320 ;
        RECT 777.470 1005.600 796.070 1465.320 ;
        RECT 799.970 1005.600 818.570 1465.320 ;
        RECT 822.470 1005.600 841.070 1465.320 ;
        RECT 844.970 1005.600 863.570 1465.320 ;
        RECT 867.470 1005.600 886.070 1465.320 ;
        RECT 889.970 1005.600 908.570 1465.320 ;
        RECT 180.615 567.820 908.570 1005.600 ;
        RECT 180.615 410.020 188.570 567.820 ;
        RECT 192.470 410.020 211.070 567.820 ;
        RECT 214.970 410.020 368.570 567.820 ;
        RECT 372.470 410.020 391.070 567.820 ;
        RECT 394.970 410.020 548.570 567.820 ;
        RECT 552.470 410.020 571.070 567.820 ;
        RECT 574.970 410.020 706.070 567.820 ;
        RECT 180.615 167.400 706.070 410.020 ;
        RECT 180.615 18.535 188.570 167.400 ;
        RECT 192.470 18.535 211.070 167.400 ;
        RECT 214.970 18.535 233.570 167.400 ;
        RECT 237.470 18.535 256.070 167.400 ;
        RECT 259.970 18.535 278.570 167.400 ;
        RECT 282.470 18.535 301.070 167.400 ;
        RECT 304.970 18.535 323.570 167.400 ;
        RECT 327.470 18.535 368.570 167.400 ;
        RECT 372.470 18.535 391.070 167.400 ;
        RECT 394.970 18.535 413.570 167.400 ;
        RECT 417.470 18.535 436.070 167.400 ;
        RECT 439.970 18.535 458.570 167.400 ;
        RECT 462.470 18.535 481.070 167.400 ;
        RECT 484.970 18.535 503.570 167.400 ;
        RECT 507.470 18.535 548.570 167.400 ;
        RECT 552.470 18.535 571.070 167.400 ;
        RECT 574.970 18.535 593.570 167.400 ;
        RECT 597.470 18.535 616.070 167.400 ;
        RECT 619.970 18.535 638.570 167.400 ;
        RECT 642.470 18.535 661.070 167.400 ;
        RECT 664.970 18.535 683.570 167.400 ;
        RECT 687.470 18.535 706.070 167.400 ;
        RECT 709.970 18.535 728.570 567.820 ;
        RECT 732.470 18.535 751.070 567.820 ;
        RECT 754.970 18.535 773.570 567.820 ;
        RECT 777.470 18.535 796.070 567.820 ;
        RECT 799.970 18.535 818.570 567.820 ;
        RECT 822.470 18.535 841.070 567.820 ;
        RECT 844.970 18.535 863.570 567.820 ;
        RECT 867.470 18.535 886.070 567.820 ;
        RECT 889.970 18.535 908.570 567.820 ;
        RECT 912.470 18.535 931.070 1465.320 ;
        RECT 934.970 18.535 953.570 3355.040 ;
        RECT 957.470 18.535 976.070 3355.040 ;
        RECT 979.970 18.535 998.570 3355.040 ;
        RECT 1002.470 18.535 1021.070 3355.040 ;
        RECT 1024.970 18.535 1043.570 3355.040 ;
        RECT 1047.470 18.535 1066.070 3355.040 ;
        RECT 1069.970 1246.850 1088.570 3355.040 ;
        RECT 1092.470 1246.850 1111.070 3355.040 ;
        RECT 1114.970 1246.850 1133.570 3355.040 ;
        RECT 1137.470 1246.850 1156.070 3355.040 ;
        RECT 1159.970 1246.850 1178.570 3355.040 ;
        RECT 1069.970 990.400 1178.570 1246.850 ;
        RECT 1069.970 18.535 1088.570 990.400 ;
        RECT 1092.470 18.535 1111.070 990.400 ;
        RECT 1114.970 18.535 1133.570 990.400 ;
        RECT 1137.470 18.535 1156.070 990.400 ;
        RECT 1159.970 18.535 1178.570 990.400 ;
        RECT 1182.470 18.535 1201.070 3355.040 ;
        RECT 1204.970 18.535 1223.570 3355.040 ;
        RECT 1227.470 18.535 1246.070 3355.040 ;
        RECT 1249.970 18.535 1268.570 3355.040 ;
        RECT 1272.470 18.535 1291.070 3355.040 ;
        RECT 1294.970 18.535 1313.570 3355.040 ;
        RECT 1317.470 18.535 1336.070 3355.040 ;
        RECT 1339.970 18.535 1358.570 3355.040 ;
        RECT 1362.470 18.535 1381.070 3355.040 ;
        RECT 1384.970 18.535 1403.570 3355.040 ;
        RECT 1407.470 18.535 1426.070 3355.040 ;
        RECT 1429.970 18.535 1448.570 3355.040 ;
        RECT 1452.470 18.535 1471.070 3355.040 ;
        RECT 1474.970 18.535 1493.570 3355.040 ;
        RECT 1497.470 18.535 1516.070 3355.040 ;
        RECT 1519.970 18.535 1538.570 3355.040 ;
        RECT 1542.470 18.535 1561.070 3355.040 ;
        RECT 1564.970 18.535 1583.570 3355.040 ;
        RECT 1587.470 613.220 1606.070 3355.040 ;
        RECT 1609.970 613.220 1628.570 3355.040 ;
        RECT 1632.470 613.220 1651.070 3355.040 ;
        RECT 1654.970 613.220 1673.570 3355.040 ;
        RECT 1677.470 3019.340 2213.570 3355.040 ;
        RECT 1677.470 2742.500 1696.070 3019.340 ;
        RECT 1699.970 2742.500 1718.570 3019.340 ;
        RECT 1722.470 2742.500 1741.070 3019.340 ;
        RECT 1744.970 2742.500 1808.570 3019.340 ;
        RECT 1812.470 2742.500 1831.070 3019.340 ;
        RECT 1834.970 2742.500 1853.570 3019.340 ;
        RECT 1857.470 2742.500 1876.070 3019.340 ;
        RECT 1879.970 2742.500 1898.570 3019.340 ;
        RECT 1902.470 2742.500 1921.070 3019.340 ;
        RECT 1924.970 2742.500 1988.570 3019.340 ;
        RECT 1992.470 2742.500 2011.070 3019.340 ;
        RECT 2014.970 2742.500 2033.570 3019.340 ;
        RECT 2037.470 2742.500 2056.070 3019.340 ;
        RECT 2059.970 2742.500 2078.570 3019.340 ;
        RECT 2082.470 2742.500 2101.070 3019.340 ;
        RECT 2104.970 2742.500 2168.570 3019.340 ;
        RECT 2172.470 2742.500 2191.070 3019.340 ;
        RECT 2194.970 2742.500 2213.570 3019.340 ;
        RECT 2217.470 2742.500 2236.070 3355.040 ;
        RECT 2239.970 2742.500 2258.570 3355.040 ;
        RECT 2262.470 2742.500 2281.070 3355.040 ;
        RECT 2284.970 2742.500 2303.570 3355.040 ;
        RECT 2307.470 2742.500 2326.070 3355.040 ;
        RECT 2329.970 2742.500 2348.570 3355.040 ;
        RECT 2352.470 2742.500 2371.070 3355.040 ;
        RECT 2374.970 2742.500 2393.570 3355.040 ;
        RECT 2397.470 2742.500 2416.070 3355.040 ;
        RECT 1677.470 2051.080 2416.070 2742.500 ;
        RECT 1677.470 1840.360 1808.570 2051.080 ;
        RECT 1812.470 1840.360 1831.070 2051.080 ;
        RECT 1834.970 1840.360 1853.570 2051.080 ;
        RECT 1857.470 1840.360 1988.570 2051.080 ;
        RECT 1992.470 1840.360 2011.070 2051.080 ;
        RECT 2014.970 1840.360 2033.570 2051.080 ;
        RECT 2037.470 1840.360 2168.570 2051.080 ;
        RECT 2172.470 1840.360 2191.070 2051.080 ;
        RECT 2194.970 1840.360 2213.570 2051.080 ;
        RECT 1677.470 1495.060 2213.570 1840.360 ;
        RECT 1677.470 1224.180 1763.570 1495.060 ;
        RECT 1767.470 1224.180 1786.070 1495.060 ;
        RECT 1789.970 1224.180 1808.570 1495.060 ;
        RECT 1812.470 1224.180 1831.070 1495.060 ;
        RECT 1834.970 1224.180 1943.570 1495.060 ;
        RECT 1947.470 1224.180 1966.070 1495.060 ;
        RECT 1969.970 1224.180 1988.570 1495.060 ;
        RECT 1992.470 1224.180 2011.070 1495.060 ;
        RECT 2014.970 1224.180 2123.570 1495.060 ;
        RECT 2127.470 1224.180 2146.070 1495.060 ;
        RECT 2149.970 1224.180 2168.570 1495.060 ;
        RECT 2172.470 1224.180 2191.070 1495.060 ;
        RECT 2194.970 1224.180 2213.570 1495.060 ;
        RECT 2217.470 1224.180 2236.070 2051.080 ;
        RECT 2239.970 1224.180 2258.570 2051.080 ;
        RECT 2262.470 1224.180 2281.070 2051.080 ;
        RECT 2284.970 1224.180 2303.570 2051.080 ;
        RECT 2307.470 1224.180 2326.070 2051.080 ;
        RECT 2329.970 1224.180 2348.570 2051.080 ;
        RECT 2352.470 1224.180 2371.070 2051.080 ;
        RECT 2374.970 1224.180 2393.570 2051.080 ;
        RECT 2397.470 1224.180 2416.070 2051.080 ;
        RECT 1677.470 786.400 2416.070 1224.180 ;
        RECT 1677.470 613.220 1808.570 786.400 ;
        RECT 1812.470 613.220 1831.070 786.400 ;
        RECT 1834.970 613.220 1988.570 786.400 ;
        RECT 1992.470 613.220 2011.070 786.400 ;
        RECT 2014.970 613.220 2123.570 786.400 ;
        RECT 1587.470 190.400 2123.570 613.220 ;
        RECT 1587.470 18.535 1606.070 190.400 ;
        RECT 1609.970 18.535 1628.570 190.400 ;
        RECT 1632.470 18.535 1651.070 190.400 ;
        RECT 1654.970 18.535 1673.570 190.400 ;
        RECT 1677.470 18.535 1696.070 190.400 ;
        RECT 1699.970 18.535 1718.570 190.400 ;
        RECT 1722.470 18.535 1741.070 190.400 ;
        RECT 1744.970 18.535 1763.570 190.400 ;
        RECT 1767.470 18.535 1786.070 190.400 ;
        RECT 1789.970 18.535 1808.570 190.400 ;
        RECT 1812.470 18.535 1831.070 190.400 ;
        RECT 1834.970 18.535 1853.570 190.400 ;
        RECT 1857.470 18.535 1876.070 190.400 ;
        RECT 1879.970 18.535 1898.570 190.400 ;
        RECT 1902.470 18.535 1921.070 190.400 ;
        RECT 1924.970 18.535 1943.570 190.400 ;
        RECT 1947.470 18.535 1966.070 190.400 ;
        RECT 1969.970 18.535 1988.570 190.400 ;
        RECT 1992.470 18.535 2011.070 190.400 ;
        RECT 2014.970 18.535 2033.570 190.400 ;
        RECT 2037.470 18.535 2056.070 190.400 ;
        RECT 2059.970 18.535 2078.570 190.400 ;
        RECT 2082.470 18.535 2101.070 190.400 ;
        RECT 2104.970 18.535 2123.570 190.400 ;
        RECT 2127.470 18.535 2146.070 786.400 ;
        RECT 2149.970 18.535 2168.570 786.400 ;
        RECT 2172.470 18.535 2191.070 786.400 ;
        RECT 2194.970 18.535 2213.570 786.400 ;
        RECT 2217.470 18.535 2236.070 786.400 ;
        RECT 2239.970 18.535 2258.570 786.400 ;
        RECT 2262.470 613.220 2348.570 786.400 ;
        RECT 2352.470 613.220 2371.070 786.400 ;
        RECT 2374.970 613.220 2416.070 786.400 ;
        RECT 2419.970 613.220 2438.570 3355.040 ;
        RECT 2442.470 613.220 2461.070 3355.040 ;
        RECT 2464.970 613.220 2483.570 3355.040 ;
        RECT 2487.470 613.220 2506.070 3355.040 ;
        RECT 2509.970 613.220 2528.570 3355.040 ;
        RECT 2532.470 613.220 2551.070 3355.040 ;
        RECT 2554.970 613.220 2573.570 3355.040 ;
        RECT 2577.470 613.220 2596.070 3355.040 ;
        RECT 2599.970 613.220 2618.570 3355.040 ;
        RECT 2622.470 613.220 2641.070 3355.040 ;
        RECT 2644.970 613.220 2663.570 3355.040 ;
        RECT 2667.470 613.220 2686.070 3355.040 ;
        RECT 2689.970 613.220 2708.570 3355.040 ;
        RECT 2712.470 613.220 2731.070 3355.040 ;
        RECT 2734.970 613.220 2753.570 3355.040 ;
        RECT 2757.470 613.220 2773.160 3355.040 ;
        RECT 2262.470 190.400 2773.160 613.220 ;
        RECT 2262.470 18.535 2281.070 190.400 ;
        RECT 2284.970 18.535 2303.570 190.400 ;
        RECT 2307.470 18.535 2326.070 190.400 ;
        RECT 2329.970 18.535 2348.570 190.400 ;
        RECT 2352.470 18.535 2371.070 190.400 ;
        RECT 2374.970 18.535 2393.570 190.400 ;
        RECT 2397.470 18.535 2416.070 190.400 ;
        RECT 2419.970 18.535 2438.570 190.400 ;
        RECT 2442.470 18.535 2461.070 190.400 ;
        RECT 2464.970 18.535 2483.570 190.400 ;
        RECT 2487.470 18.535 2506.070 190.400 ;
        RECT 2509.970 18.535 2528.570 190.400 ;
        RECT 2532.470 18.535 2551.070 190.400 ;
        RECT 2554.970 18.535 2573.570 190.400 ;
        RECT 2577.470 18.535 2596.070 190.400 ;
        RECT 2599.970 18.535 2618.570 190.400 ;
        RECT 2622.470 18.535 2641.070 190.400 ;
        RECT 2644.970 18.535 2663.570 190.400 ;
        RECT 2667.470 18.535 2686.070 190.400 ;
        RECT 2689.970 18.535 2708.570 190.400 ;
        RECT 2712.470 18.535 2731.070 190.400 ;
        RECT 2734.970 18.535 2753.570 190.400 ;
        RECT 2757.470 18.535 2773.160 190.400 ;
  END
END user_project_wrapper
END LIBRARY

